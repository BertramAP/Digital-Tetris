module Memory(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_1(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_2(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_2.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_3(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_3.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_4(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_4.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_5(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_5.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_6(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_6.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_7(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_7.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_8(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_8.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_9(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_9.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_10(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_10.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_11(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_11.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_12(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_12.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_13(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_13.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_14(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_14.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_15(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_15.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_16(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_16.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_17(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_17.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_18(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_18.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_19(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_19.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_20(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_20.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_21(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_21.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_22(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_22.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_23(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_23.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_24(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_24.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_25(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_25.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_26(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_26.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_27(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_27.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_28(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_28.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_29(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_29.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_30(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_30.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_31(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_31.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_32(
  input         clock,
  input  [10:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [4:0]  io_dataRead, // @[\\src\\main\\scala\\Memory.scala 48:14]
  input         io_writeEnable, // @[\\src\\main\\scala\\Memory.scala 48:14]
  input  [4:0]  io_dataWrite // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [10:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [4:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 57:26]
  wire [4:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 57:26]
  RamSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5)) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 57:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 63:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 58:21]
  assign ramsSpWf_we = io_writeEnable; // @[\\src\\main\\scala\\Memory.scala 59:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 60:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 61:22]
  assign ramsSpWf_di = io_dataWrite; // @[\\src\\main\\scala\\Memory.scala 62:20]
endmodule
module Memory_34(
  input         clock,
  input  [10:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [4:0]  io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [10:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [4:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [4:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5), .LOAD_FILE("memory_init/backbuffer_init.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 5'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_35(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_36(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_37(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_2.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_38(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_3.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_39(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_4.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_40(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_5.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_41(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_6.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_42(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_7.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_43(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_8.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_44(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_9.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_45(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_10.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_46(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_11.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_47(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_12.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_48(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_13.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_49(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_14.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_50(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_15.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_51(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_16.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_52(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_17.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_53(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_18.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_54(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_19.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_55(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_20.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_56(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_21.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_57(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_22.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_58(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_23.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_59(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_24.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_60(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_25.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_61(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_26.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_62(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_27.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_63(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_28.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_64(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_29.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_65(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_30.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_66(
  input        clock,
  input  [9:0] io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [6:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [9:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [6:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_31.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 7'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module MultiHotPriortyReductionTree(
  input  [5:0] io_dataInput_0, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_1, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_2, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_3, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_4, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_5, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_6, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_7, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_8, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_9, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_10, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_11, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_12, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_13, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_14, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_15, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_16, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_17, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_18, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_19, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_20, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_21, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_22, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_23, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_24, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_25, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_26, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_27, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_28, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_29, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_30, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input  [5:0] io_dataInput_31, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_0, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_1, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_2, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_3, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_4, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_5, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_6, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_7, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_8, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_9, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_10, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_11, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_12, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_13, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_14, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_15, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_16, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_17, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_18, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_19, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_20, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_21, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_22, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_23, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_24, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_25, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_26, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_27, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_28, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_29, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_30, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  input        io_selectInput_31, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  output [5:0] io_dataOutput, // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
  output       io_selectOutput // @[\\src\\main\\scala\\GameUtilities.scala 53:14]
);
  wire  selectNodeOutputs_15 = io_selectInput_0 | io_selectInput_1; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_16 = io_selectInput_2 | io_selectInput_3; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_7 = selectNodeOutputs_15 | selectNodeOutputs_16; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_17 = io_selectInput_4 | io_selectInput_5; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_18 = io_selectInput_6 | io_selectInput_7; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_8 = selectNodeOutputs_17 | selectNodeOutputs_18; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_3 = selectNodeOutputs_7 | selectNodeOutputs_8; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_19 = io_selectInput_8 | io_selectInput_9; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_20 = io_selectInput_10 | io_selectInput_11; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_9 = selectNodeOutputs_19 | selectNodeOutputs_20; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_21 = io_selectInput_12 | io_selectInput_13; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_22 = io_selectInput_14 | io_selectInput_15; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_10 = selectNodeOutputs_21 | selectNodeOutputs_22; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_4 = selectNodeOutputs_9 | selectNodeOutputs_10; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_1 = selectNodeOutputs_3 | selectNodeOutputs_4; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_15 = io_selectInput_0 ? io_dataInput_0 : io_dataInput_1; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_16 = io_selectInput_2 ? io_dataInput_2 : io_dataInput_3; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_7 = selectNodeOutputs_15 ? dataNodeOutputs_15 : dataNodeOutputs_16; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_17 = io_selectInput_4 ? io_dataInput_4 : io_dataInput_5; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_18 = io_selectInput_6 ? io_dataInput_6 : io_dataInput_7; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_8 = selectNodeOutputs_17 ? dataNodeOutputs_17 : dataNodeOutputs_18; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_3 = selectNodeOutputs_7 ? dataNodeOutputs_7 : dataNodeOutputs_8; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_19 = io_selectInput_8 ? io_dataInput_8 : io_dataInput_9; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_20 = io_selectInput_10 ? io_dataInput_10 : io_dataInput_11; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_9 = selectNodeOutputs_19 ? dataNodeOutputs_19 : dataNodeOutputs_20; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_21 = io_selectInput_12 ? io_dataInput_12 : io_dataInput_13; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_22 = io_selectInput_14 ? io_dataInput_14 : io_dataInput_15; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_10 = selectNodeOutputs_21 ? dataNodeOutputs_21 : dataNodeOutputs_22; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_4 = selectNodeOutputs_9 ? dataNodeOutputs_9 : dataNodeOutputs_10; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_1 = selectNodeOutputs_3 ? dataNodeOutputs_3 : dataNodeOutputs_4; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_23 = io_selectInput_16 | io_selectInput_17; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_24 = io_selectInput_18 | io_selectInput_19; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_11 = selectNodeOutputs_23 | selectNodeOutputs_24; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_25 = io_selectInput_20 | io_selectInput_21; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_26 = io_selectInput_22 | io_selectInput_23; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_12 = selectNodeOutputs_25 | selectNodeOutputs_26; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_5 = selectNodeOutputs_11 | selectNodeOutputs_12; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_23 = io_selectInput_16 ? io_dataInput_16 : io_dataInput_17; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_24 = io_selectInput_18 ? io_dataInput_18 : io_dataInput_19; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_11 = selectNodeOutputs_23 ? dataNodeOutputs_23 : dataNodeOutputs_24; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_25 = io_selectInput_20 ? io_dataInput_20 : io_dataInput_21; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_26 = io_selectInput_22 ? io_dataInput_22 : io_dataInput_23; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_12 = selectNodeOutputs_25 ? dataNodeOutputs_25 : dataNodeOutputs_26; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_5 = selectNodeOutputs_11 ? dataNodeOutputs_11 : dataNodeOutputs_12; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_27 = io_selectInput_24 | io_selectInput_25; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_28 = io_selectInput_26 | io_selectInput_27; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_13 = selectNodeOutputs_27 | selectNodeOutputs_28; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_27 = io_selectInput_24 ? io_dataInput_24 : io_dataInput_25; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_28 = io_selectInput_26 ? io_dataInput_26 : io_dataInput_27; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_13 = selectNodeOutputs_27 ? dataNodeOutputs_27 : dataNodeOutputs_28; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_29 = io_selectInput_28 | io_selectInput_29; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_29 = io_selectInput_28 ? io_dataInput_28 : io_dataInput_29; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_30 = io_selectInput_30 ? io_dataInput_30 : io_dataInput_31; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_14 = selectNodeOutputs_29 ? dataNodeOutputs_29 : dataNodeOutputs_30; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_6 = selectNodeOutputs_13 ? dataNodeOutputs_13 : dataNodeOutputs_14; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_2 = selectNodeOutputs_5 ? dataNodeOutputs_5 : dataNodeOutputs_6; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  wire  selectNodeOutputs_30 = io_selectInput_30 | io_selectInput_31; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_14 = selectNodeOutputs_29 | selectNodeOutputs_30; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_6 = selectNodeOutputs_13 | selectNodeOutputs_14; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  wire  selectNodeOutputs_2 = selectNodeOutputs_5 | selectNodeOutputs_6; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
  assign io_dataOutput = selectNodeOutputs_1 ? dataNodeOutputs_1 : dataNodeOutputs_2; // @[\\src\\main\\scala\\GameUtilities.scala 85:34]
  assign io_selectOutput = selectNodeOutputs_1 | selectNodeOutputs_2; // @[\\src\\main\\scala\\GameUtilities.scala 86:54]
endmodule
module GraphicEngineVGA(
  input         clock,
  input         reset,
  input  [10:0] io_spriteXPosition_0, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_1, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_2, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_4, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_5, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_6, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_15, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_spriteXPosition_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_0, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_1, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_2, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_4, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_5, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_6, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_15, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_spriteYPosition_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_0, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_1, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_2, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_3, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_4, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_5, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_6, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_7, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_8, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_9, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_10, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_11, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_12, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_13, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_14, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_15, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_16, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_17, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_18, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_19, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_20, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_21, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_22, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_23, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_24, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_25, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_26, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_spriteVisible_27, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [9:0]  io_viewBoxX, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [8:0]  io_viewBoxY, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [4:0]  io_backBufferWriteData, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input  [10:0] io_backBufferWriteAddress, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_backBufferWriteEnable, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_newFrame, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  input         io_frameUpdateDone, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_missingFrameError, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_backBufferWriteError, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_viewBoxOutOfRangeError, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaRed, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaBlue, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output [3:0]  io_vgaGreen, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_Hsync, // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
  output        io_Vsync // @[\\src\\main\\scala\\GraphicEngineVGA.scala 12:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
`endif // RANDOMIZE_REG_INIT
  wire  backTileMemories_0_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_0_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_1_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_1_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_2_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_2_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_3_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_3_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_4_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_4_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_5_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_5_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_6_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_6_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_7_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_7_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_8_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_8_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_9_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_9_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_10_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_10_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_11_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_11_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_12_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_12_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_13_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_13_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_14_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_14_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_15_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_15_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_16_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_16_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_17_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_17_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_18_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_18_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_19_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_19_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_20_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_20_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_21_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_21_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_22_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_22_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_23_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_23_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_24_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_24_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_25_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_25_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_26_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_26_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_27_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_27_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_28_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_28_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_29_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_29_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_30_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_30_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backTileMemories_31_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [9:0] backTileMemories_31_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire [6:0] backTileMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
  wire  backBufferMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [10:0] backBufferMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [4:0] backBufferMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire  backBufferMemory_io_writeEnable; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire [4:0] backBufferMemory_io_dataWrite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
  wire  backBufferShadowMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [10:0] backBufferShadowMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [4:0] backBufferShadowMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire  backBufferShadowMemory_io_writeEnable; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire [4:0] backBufferShadowMemory_io_dataWrite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
  wire  backBufferRestoreMemory_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire [10:0] backBufferRestoreMemory_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire [4:0] backBufferRestoreMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
  wire  spriteMemories_0_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_0_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_1_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_1_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_2_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_2_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_3_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_3_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_4_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_4_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_5_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_5_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_6_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_6_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_7_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_7_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_8_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_8_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_9_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_9_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_10_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_10_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_11_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_11_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_12_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_12_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_13_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_13_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_14_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_14_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_15_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_15_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_16_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_16_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_17_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_17_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_18_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_18_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_19_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_19_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_20_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_20_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_21_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_21_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_22_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_22_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_23_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_23_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_24_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_24_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_25_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_25_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_26_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_26_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_27_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_27_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_28_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_28_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_29_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_29_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_30_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_30_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire  spriteMemories_31_clock; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [9:0] spriteMemories_31_io_address; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [6:0] spriteMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectInput_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  wire  multiHotPriortyReductionTree_io_selectOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
  reg [1:0] ScaleCounterReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
  reg [9:0] CounterXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
  reg [9:0] CounterYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
  wire  _T_2 = CounterYReg == 10'h20c; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 78:26]
  wire [9:0] _CounterYReg_T_1 = CounterYReg + 10'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 82:38]
  wire [9:0] _GEN_0 = CounterYReg == 10'h20c ? 10'h0 : _CounterYReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 78:131 79:23 82:23]
  wire [9:0] _CounterXReg_T_1 = CounterXReg + 10'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 85:36]
  wire  _GEN_4 = CounterXReg == 10'h31f & _T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129 71:15]
  wire [1:0] _ScaleCounterReg_T_1 = ScaleCounterReg + 2'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 88:42]
  wire  _GEN_8 = ScaleCounterReg == 2'h3 & _GEN_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 71:15 74:52]
  reg [11:0] backMemoryRestoreCounter; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
  wire  restoreEnabled = backMemoryRestoreCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:33]
  wire  run = restoreEnabled ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:70 209:9 213:9]
  wire  Hsync = CounterXReg >= 10'h290 & CounterXReg < 10'h2f0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 92:79]
  wire  Vsync = CounterYReg >= 10'h1ea & CounterYReg < 10'h1ec; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 93:79]
  reg  io_Hsync_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Hsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  io_Vsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg [20:0] frameClockCount; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
  wire [20:0] _frameClockCount_T_2 = frameClockCount + 21'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 105:92]
  wire  preDisplayArea = frameClockCount >= 21'h199a1b; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 106:40]
  reg [10:0] spriteXPositionReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [10:0] spriteXPositionReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
  reg [9:0] spriteYPositionReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg [9:0] spriteYPositionReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
  reg  spriteVisibleReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  reg  spriteVisibleReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:35]
  wire  _GEN_77 = io_newFrame ? io_spriteVisible_0 : spriteVisibleReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_78 = io_newFrame ? io_spriteVisible_1 : spriteVisibleReg_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_79 = io_newFrame ? io_spriteVisible_2 : spriteVisibleReg_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_80 = io_newFrame ? io_spriteVisible_3 : spriteVisibleReg_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_81 = io_newFrame ? io_spriteVisible_4 : spriteVisibleReg_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_82 = io_newFrame ? io_spriteVisible_5 : spriteVisibleReg_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_83 = io_newFrame ? io_spriteVisible_6 : spriteVisibleReg_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_84 = io_newFrame ? io_spriteVisible_7 : spriteVisibleReg_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_85 = io_newFrame ? io_spriteVisible_8 : spriteVisibleReg_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_86 = io_newFrame ? io_spriteVisible_9 : spriteVisibleReg_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_87 = io_newFrame ? io_spriteVisible_10 : spriteVisibleReg_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_88 = io_newFrame ? io_spriteVisible_11 : spriteVisibleReg_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_89 = io_newFrame ? io_spriteVisible_12 : spriteVisibleReg_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_90 = io_newFrame ? io_spriteVisible_13 : spriteVisibleReg_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_91 = io_newFrame ? io_spriteVisible_14 : spriteVisibleReg_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_92 = io_newFrame ? io_spriteVisible_15 : spriteVisibleReg_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_93 = io_newFrame ? io_spriteVisible_16 : spriteVisibleReg_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_94 = io_newFrame ? io_spriteVisible_17 : spriteVisibleReg_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_95 = io_newFrame ? io_spriteVisible_18 : spriteVisibleReg_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_96 = io_newFrame ? io_spriteVisible_19 : spriteVisibleReg_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_97 = io_newFrame ? io_spriteVisible_20 : spriteVisibleReg_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_98 = io_newFrame ? io_spriteVisible_21 : spriteVisibleReg_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_99 = io_newFrame ? io_spriteVisible_22 : spriteVisibleReg_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_100 = io_newFrame ? io_spriteVisible_23 : spriteVisibleReg_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_101 = io_newFrame ? io_spriteVisible_24 : spriteVisibleReg_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_102 = io_newFrame ? io_spriteVisible_25 : spriteVisibleReg_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_103 = io_newFrame ? io_spriteVisible_26 : spriteVisibleReg_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_104 = io_newFrame ? io_spriteVisible_27 : spriteVisibleReg_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_105 = io_newFrame ? 1'h0 : spriteVisibleReg_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_106 = io_newFrame ? 1'h0 : spriteVisibleReg_29; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_107 = io_newFrame ? 1'h0 : spriteVisibleReg_30; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  wire  _GEN_108 = io_newFrame ? 1'h0 : spriteVisibleReg_31; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35,35}]
  reg [9:0] viewBoxXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
  reg [8:0] viewBoxYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
  reg  missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
  reg  backBufferWriteErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 129:40]
  reg  viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
  wire [9:0] viewBoxXClipped = viewBoxXReg >= 10'h280 ? 10'h280 : viewBoxXReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 137:28]
  wire [8:0] viewBoxYClipped = viewBoxYReg >= 9'h1e0 ? 9'h1e0 : viewBoxYReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 138:28]
  wire [10:0] pixelXBack = CounterXReg + viewBoxXClipped; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 139:27]
  wire [9:0] _GEN_860 = {{1'd0}, viewBoxYClipped}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 140:27]
  wire [10:0] pixelYBack = CounterYReg + _GEN_860; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 140:27]
  wire  _GEN_303 = viewBoxXReg > 10'h280 | viewBoxYReg > 9'h1e0 | viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 141:51 142:31 130:42]
  reg  newFrameStikyReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
  wire  _GEN_304 = io_newFrame | newFrameStikyReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 148:21 149:22 147:33]
  reg  REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:16]
  wire  _GEN_306 = newFrameStikyReg & io_newFrame | missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 154:41 155:26 128:37]
  wire [10:0] _backTileMemories_0_io_address_T_2 = 6'h20 * pixelYBack[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:75]
  wire [10:0] _GEN_861 = {{6'd0}, pixelXBack[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:62]
  wire [11:0] _backTileMemories_0_io_address_T_3 = _GEN_861 + _backTileMemories_0_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:62]
  reg [6:0] backTileMemoryDataRead_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [6:0] backTileMemoryDataRead_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
  reg [11:0] backMemoryCopyCounter; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
  wire  _T_7 = backMemoryCopyCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 187:32]
  wire [11:0] _backMemoryCopyCounter_T_1 = backMemoryCopyCounter + 12'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 188:54]
  wire  copyEnabled = preDisplayArea & _T_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23 198:17]
  reg  copyEnabledReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 200:31]
  wire [11:0] _backMemoryRestoreCounter_T_1 = backMemoryRestoreCounter + 12'h1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 206:58]
  reg [10:0] backBufferShadowMemory_io_address_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:67]
  reg [10:0] backBufferShadowMemory_io_address_REG_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:156]
  wire [10:0] _backBufferShadowMemory_io_address_T_2 = copyEnabled ? backMemoryCopyCounter[10:0] :
    backBufferShadowMemory_io_address_REG_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:105]
  reg  backBufferShadowMemory_io_writeEnable_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:71]
  reg  backBufferShadowMemory_io_writeEnable_REG_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:122]
  wire  _backBufferShadowMemory_io_writeEnable_T = copyEnabled ? 1'h0 : backBufferShadowMemory_io_writeEnable_REG_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:92]
  reg [4:0] backBufferShadowMemory_io_dataWrite_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 224:106]
  reg [10:0] backBufferMemory_io_address_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:61]
  wire [11:0] _backBufferMemory_io_address_T_3 = 6'h28 * pixelYBack[10:5]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:130]
  wire [11:0] _GEN_893 = {{6'd0}, pixelXBack[10:5]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:117]
  wire [12:0] _backBufferMemory_io_address_T_4 = _GEN_893 + _backBufferMemory_io_address_T_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:117]
  wire [12:0] _backBufferMemory_io_address_T_5 = copyEnabledReg ? {{2'd0}, backBufferMemory_io_address_REG} :
    _backBufferMemory_io_address_T_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:37]
  wire  _GEN_314 = io_backBufferWriteEnable | backBufferWriteErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 234:36 235:31 129:40]
  reg [4:0] fullBackgroundColor_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:56]
  wire [6:0] _GEN_317 = 5'h1 == fullBackgroundColor_REG ? backTileMemoryDataRead_1_REG : backTileMemoryDataRead_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_318 = 5'h2 == fullBackgroundColor_REG ? backTileMemoryDataRead_2_REG : _GEN_317; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_319 = 5'h3 == fullBackgroundColor_REG ? backTileMemoryDataRead_3_REG : _GEN_318; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_320 = 5'h4 == fullBackgroundColor_REG ? backTileMemoryDataRead_4_REG : _GEN_319; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_321 = 5'h5 == fullBackgroundColor_REG ? backTileMemoryDataRead_5_REG : _GEN_320; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_322 = 5'h6 == fullBackgroundColor_REG ? backTileMemoryDataRead_6_REG : _GEN_321; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_323 = 5'h7 == fullBackgroundColor_REG ? backTileMemoryDataRead_7_REG : _GEN_322; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_324 = 5'h8 == fullBackgroundColor_REG ? backTileMemoryDataRead_8_REG : _GEN_323; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_325 = 5'h9 == fullBackgroundColor_REG ? backTileMemoryDataRead_9_REG : _GEN_324; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_326 = 5'ha == fullBackgroundColor_REG ? backTileMemoryDataRead_10_REG : _GEN_325; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_327 = 5'hb == fullBackgroundColor_REG ? backTileMemoryDataRead_11_REG : _GEN_326; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_328 = 5'hc == fullBackgroundColor_REG ? backTileMemoryDataRead_12_REG : _GEN_327; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_329 = 5'hd == fullBackgroundColor_REG ? backTileMemoryDataRead_13_REG : _GEN_328; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_330 = 5'he == fullBackgroundColor_REG ? backTileMemoryDataRead_14_REG : _GEN_329; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_331 = 5'hf == fullBackgroundColor_REG ? backTileMemoryDataRead_15_REG : _GEN_330; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_332 = 5'h10 == fullBackgroundColor_REG ? backTileMemoryDataRead_16_REG : _GEN_331; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_333 = 5'h11 == fullBackgroundColor_REG ? backTileMemoryDataRead_17_REG : _GEN_332; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_334 = 5'h12 == fullBackgroundColor_REG ? backTileMemoryDataRead_18_REG : _GEN_333; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_335 = 5'h13 == fullBackgroundColor_REG ? backTileMemoryDataRead_19_REG : _GEN_334; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_336 = 5'h14 == fullBackgroundColor_REG ? backTileMemoryDataRead_20_REG : _GEN_335; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_337 = 5'h15 == fullBackgroundColor_REG ? backTileMemoryDataRead_21_REG : _GEN_336; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_338 = 5'h16 == fullBackgroundColor_REG ? backTileMemoryDataRead_22_REG : _GEN_337; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_339 = 5'h17 == fullBackgroundColor_REG ? backTileMemoryDataRead_23_REG : _GEN_338; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_340 = 5'h18 == fullBackgroundColor_REG ? backTileMemoryDataRead_24_REG : _GEN_339; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_341 = 5'h19 == fullBackgroundColor_REG ? backTileMemoryDataRead_25_REG : _GEN_340; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_342 = 5'h1a == fullBackgroundColor_REG ? backTileMemoryDataRead_26_REG : _GEN_341; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_343 = 5'h1b == fullBackgroundColor_REG ? backTileMemoryDataRead_27_REG : _GEN_342; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_344 = 5'h1c == fullBackgroundColor_REG ? backTileMemoryDataRead_28_REG : _GEN_343; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_345 = 5'h1d == fullBackgroundColor_REG ? backTileMemoryDataRead_29_REG : _GEN_344; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] _GEN_346 = 5'h1e == fullBackgroundColor_REG ? backTileMemoryDataRead_30_REG : _GEN_345; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  wire [6:0] fullBackgroundColor = 5'h1f == fullBackgroundColor_REG ? backTileMemoryDataRead_31_REG : _GEN_346; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:{23,23}]
  reg [5:0] pixelColorBack; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 245:31]
  wire [10:0] _inSpriteXValue_T_1 = {1'h0,CounterXReg}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:47]
  wire [11:0] inSpriteXValue = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_0); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_0 = $signed(inSpriteXValue) >= 12'sh0 & $signed(inSpriteXValue) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_354 = {{1{inSpriteXValue[11]}},inSpriteXValue}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _inSpriteYValue_T_1 = {1'h0,CounterYReg}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:47]
  wire [10:0] _GEN_894 = {{1{spriteYPositionReg_0[9]}},spriteYPositionReg_0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue = $signed(_inSpriteYValue_T_1) - $signed(_GEN_894); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_0 = inSpriteYValue[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_0 = $signed(inSpriteYPreScaled_0) >= 11'sh0 & $signed(inSpriteYPreScaled_0) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_362 = {{1{inSpriteYPreScaled_0[10]}},inSpriteYPreScaled_0}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_1 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_1); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_1 = $signed(inSpriteXValue_1) >= 12'sh0 & $signed(inSpriteXValue_1) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_370 = {{1{inSpriteXValue_1[11]}},inSpriteXValue_1}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_896 = {{1{spriteYPositionReg_1[9]}},spriteYPositionReg_1}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_1 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_896); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_1 = inSpriteYValue_1[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_1 = $signed(inSpriteYPreScaled_1) >= 11'sh0 & $signed(inSpriteYPreScaled_1) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_378 = {{1{inSpriteYPreScaled_1[10]}},inSpriteYPreScaled_1}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_2 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_2); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_2 = $signed(inSpriteXValue_2) >= 12'sh0 & $signed(inSpriteXValue_2) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_386 = {{1{inSpriteXValue_2[11]}},inSpriteXValue_2}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_898 = {{1{spriteYPositionReg_2[9]}},spriteYPositionReg_2}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_2 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_898); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_2 = inSpriteYValue_2[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_2 = $signed(inSpriteYPreScaled_2) >= 11'sh0 & $signed(inSpriteYPreScaled_2) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_394 = {{1{inSpriteYPreScaled_2[10]}},inSpriteYPreScaled_2}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_3 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_3); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_3 = $signed(inSpriteXValue_3) >= 12'sh0 & $signed(inSpriteXValue_3) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_402 = {{1{inSpriteXValue_3[11]}},inSpriteXValue_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_900 = {{1{spriteYPositionReg_3[9]}},spriteYPositionReg_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_3 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_900); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_3 = inSpriteYValue_3[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_3 = $signed(inSpriteYPreScaled_3) >= 11'sh0 & $signed(inSpriteYPreScaled_3) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_410 = {{1{inSpriteYPreScaled_3[10]}},inSpriteYPreScaled_3}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_4 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_4); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_4 = $signed(inSpriteXValue_4) >= 12'sh0 & $signed(inSpriteXValue_4) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_418 = {{1{inSpriteXValue_4[11]}},inSpriteXValue_4}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_902 = {{1{spriteYPositionReg_4[9]}},spriteYPositionReg_4}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_4 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_902); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_4 = inSpriteYValue_4[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_4 = $signed(inSpriteYPreScaled_4) >= 11'sh0 & $signed(inSpriteYPreScaled_4) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_426 = {{1{inSpriteYPreScaled_4[10]}},inSpriteYPreScaled_4}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_5 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_5); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_5 = $signed(inSpriteXValue_5) >= 12'sh0 & $signed(inSpriteXValue_5) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_434 = {{1{inSpriteXValue_5[11]}},inSpriteXValue_5}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_904 = {{1{spriteYPositionReg_5[9]}},spriteYPositionReg_5}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_5 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_904); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_5 = inSpriteYValue_5[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_5 = $signed(inSpriteYPreScaled_5) >= 11'sh0 & $signed(inSpriteYPreScaled_5) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_442 = {{1{inSpriteYPreScaled_5[10]}},inSpriteYPreScaled_5}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_6 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_6); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_6 = $signed(inSpriteXValue_6) >= 12'sh0 & $signed(inSpriteXValue_6) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_450 = {{1{inSpriteXValue_6[11]}},inSpriteXValue_6}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_906 = {{1{spriteYPositionReg_6[9]}},spriteYPositionReg_6}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_6 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_906); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_6 = inSpriteYValue_6[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_6 = $signed(inSpriteYPreScaled_6) >= 11'sh0 & $signed(inSpriteYPreScaled_6) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_458 = {{1{inSpriteYPreScaled_6[10]}},inSpriteYPreScaled_6}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_7 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_7); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_7 = $signed(inSpriteXValue_7) >= 12'sh0 & $signed(inSpriteXValue_7) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_466 = {{1{inSpriteXValue_7[11]}},inSpriteXValue_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_908 = {{1{spriteYPositionReg_7[9]}},spriteYPositionReg_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_7 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_908); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_7 = inSpriteYValue_7[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_7 = $signed(inSpriteYPreScaled_7) >= 11'sh0 & $signed(inSpriteYPreScaled_7) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_474 = {{1{inSpriteYPreScaled_7[10]}},inSpriteYPreScaled_7}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_8 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_8); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_8 = $signed(inSpriteXValue_8) >= 12'sh0 & $signed(inSpriteXValue_8) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_482 = {{1{inSpriteXValue_8[11]}},inSpriteXValue_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_910 = {{1{spriteYPositionReg_8[9]}},spriteYPositionReg_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_8 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_910); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_8 = inSpriteYValue_8[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_8 = $signed(inSpriteYPreScaled_8) >= 11'sh0 & $signed(inSpriteYPreScaled_8) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_490 = {{1{inSpriteYPreScaled_8[10]}},inSpriteYPreScaled_8}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_9 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_9); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_9 = $signed(inSpriteXValue_9) >= 12'sh0 & $signed(inSpriteXValue_9) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_498 = {{1{inSpriteXValue_9[11]}},inSpriteXValue_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_912 = {{1{spriteYPositionReg_9[9]}},spriteYPositionReg_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_9 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_912); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_9 = inSpriteYValue_9[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_9 = $signed(inSpriteYPreScaled_9) >= 11'sh0 & $signed(inSpriteYPreScaled_9) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_506 = {{1{inSpriteYPreScaled_9[10]}},inSpriteYPreScaled_9}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_10 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_10); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_10 = $signed(inSpriteXValue_10) >= 12'sh0 & $signed(inSpriteXValue_10) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_514 = {{1{inSpriteXValue_10[11]}},inSpriteXValue_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_914 = {{1{spriteYPositionReg_10[9]}},spriteYPositionReg_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_10 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_914); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_10 = inSpriteYValue_10[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_10 = $signed(inSpriteYPreScaled_10) >= 11'sh0 & $signed(inSpriteYPreScaled_10) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_522 = {{1{inSpriteYPreScaled_10[10]}},inSpriteYPreScaled_10}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_11 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_11); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_11 = $signed(inSpriteXValue_11) >= 12'sh0 & $signed(inSpriteXValue_11) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_530 = {{1{inSpriteXValue_11[11]}},inSpriteXValue_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_916 = {{1{spriteYPositionReg_11[9]}},spriteYPositionReg_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_11 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_916); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_11 = inSpriteYValue_11[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_11 = $signed(inSpriteYPreScaled_11) >= 11'sh0 & $signed(inSpriteYPreScaled_11) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_538 = {{1{inSpriteYPreScaled_11[10]}},inSpriteYPreScaled_11}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_12 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_12); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_12 = $signed(inSpriteXValue_12) >= 12'sh0 & $signed(inSpriteXValue_12) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_546 = {{1{inSpriteXValue_12[11]}},inSpriteXValue_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_918 = {{1{spriteYPositionReg_12[9]}},spriteYPositionReg_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_12 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_918); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_12 = inSpriteYValue_12[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_12 = $signed(inSpriteYPreScaled_12) >= 11'sh0 & $signed(inSpriteYPreScaled_12) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_554 = {{1{inSpriteYPreScaled_12[10]}},inSpriteYPreScaled_12}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_13 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_13); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_13 = $signed(inSpriteXValue_13) >= 12'sh0 & $signed(inSpriteXValue_13) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_562 = {{1{inSpriteXValue_13[11]}},inSpriteXValue_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_920 = {{1{spriteYPositionReg_13[9]}},spriteYPositionReg_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_13 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_920); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_13 = inSpriteYValue_13[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_13 = $signed(inSpriteYPreScaled_13) >= 11'sh0 & $signed(inSpriteYPreScaled_13) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_570 = {{1{inSpriteYPreScaled_13[10]}},inSpriteYPreScaled_13}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_14 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_14); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_14 = $signed(inSpriteXValue_14) >= 12'sh0 & $signed(inSpriteXValue_14) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_578 = {{1{inSpriteXValue_14[11]}},inSpriteXValue_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_922 = {{1{spriteYPositionReg_14[9]}},spriteYPositionReg_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_14 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_922); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_14 = inSpriteYValue_14[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_14 = $signed(inSpriteYPreScaled_14) >= 11'sh0 & $signed(inSpriteYPreScaled_14) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_586 = {{1{inSpriteYPreScaled_14[10]}},inSpriteYPreScaled_14}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_15 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_15); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_15 = $signed(inSpriteXValue_15) >= 12'sh0 & $signed(inSpriteXValue_15) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_594 = {{1{inSpriteXValue_15[11]}},inSpriteXValue_15}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_924 = {{1{spriteYPositionReg_15[9]}},spriteYPositionReg_15}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_15 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_924); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_15 = inSpriteYValue_15[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_15 = $signed(inSpriteYPreScaled_15) >= 11'sh0 & $signed(inSpriteYPreScaled_15) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_602 = {{1{inSpriteYPreScaled_15[10]}},inSpriteYPreScaled_15}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_16 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_16); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_16 = $signed(inSpriteXValue_16) >= 12'sh0 & $signed(inSpriteXValue_16) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_610 = {{1{inSpriteXValue_16[11]}},inSpriteXValue_16}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_926 = {{1{spriteYPositionReg_16[9]}},spriteYPositionReg_16}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_16 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_926); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_16 = inSpriteYValue_16[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_16 = $signed(inSpriteYPreScaled_16) >= 11'sh0 & $signed(inSpriteYPreScaled_16) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_618 = {{1{inSpriteYPreScaled_16[10]}},inSpriteYPreScaled_16}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_17 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_17); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_17 = $signed(inSpriteXValue_17) >= 12'sh0 & $signed(inSpriteXValue_17) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_626 = {{1{inSpriteXValue_17[11]}},inSpriteXValue_17}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_928 = {{1{spriteYPositionReg_17[9]}},spriteYPositionReg_17}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_17 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_928); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_17 = inSpriteYValue_17[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_17 = $signed(inSpriteYPreScaled_17) >= 11'sh0 & $signed(inSpriteYPreScaled_17) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_634 = {{1{inSpriteYPreScaled_17[10]}},inSpriteYPreScaled_17}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_18 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_18); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_18 = $signed(inSpriteXValue_18) >= 12'sh0 & $signed(inSpriteXValue_18) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_642 = {{1{inSpriteXValue_18[11]}},inSpriteXValue_18}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_930 = {{1{spriteYPositionReg_18[9]}},spriteYPositionReg_18}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_18 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_930); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_18 = inSpriteYValue_18[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_18 = $signed(inSpriteYPreScaled_18) >= 11'sh0 & $signed(inSpriteYPreScaled_18) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_650 = {{1{inSpriteYPreScaled_18[10]}},inSpriteYPreScaled_18}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_19 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_19); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_19 = $signed(inSpriteXValue_19) >= 12'sh0 & $signed(inSpriteXValue_19) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_658 = {{1{inSpriteXValue_19[11]}},inSpriteXValue_19}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_932 = {{1{spriteYPositionReg_19[9]}},spriteYPositionReg_19}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_19 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_932); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_19 = inSpriteYValue_19[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_19 = $signed(inSpriteYPreScaled_19) >= 11'sh0 & $signed(inSpriteYPreScaled_19) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_666 = {{1{inSpriteYPreScaled_19[10]}},inSpriteYPreScaled_19}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_20 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_20); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_20 = $signed(inSpriteXValue_20) >= 12'sh0 & $signed(inSpriteXValue_20) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_674 = {{1{inSpriteXValue_20[11]}},inSpriteXValue_20}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_934 = {{1{spriteYPositionReg_20[9]}},spriteYPositionReg_20}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_20 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_934); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_20 = inSpriteYValue_20[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_20 = $signed(inSpriteYPreScaled_20) >= 11'sh0 & $signed(inSpriteYPreScaled_20) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_682 = {{1{inSpriteYPreScaled_20[10]}},inSpriteYPreScaled_20}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_21 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_21); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_21 = $signed(inSpriteXValue_21) >= 12'sh0 & $signed(inSpriteXValue_21) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_690 = {{1{inSpriteXValue_21[11]}},inSpriteXValue_21}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_936 = {{1{spriteYPositionReg_21[9]}},spriteYPositionReg_21}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_21 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_936); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_21 = inSpriteYValue_21[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_21 = $signed(inSpriteYPreScaled_21) >= 11'sh0 & $signed(inSpriteYPreScaled_21) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_698 = {{1{inSpriteYPreScaled_21[10]}},inSpriteYPreScaled_21}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_22 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_22); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_22 = $signed(inSpriteXValue_22) >= 12'sh0 & $signed(inSpriteXValue_22) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_706 = {{1{inSpriteXValue_22[11]}},inSpriteXValue_22}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_938 = {{1{spriteYPositionReg_22[9]}},spriteYPositionReg_22}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_22 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_938); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_22 = inSpriteYValue_22[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_22 = $signed(inSpriteYPreScaled_22) >= 11'sh0 & $signed(inSpriteYPreScaled_22) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_714 = {{1{inSpriteYPreScaled_22[10]}},inSpriteYPreScaled_22}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_23 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_23); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_23 = $signed(inSpriteXValue_23) >= 12'sh0 & $signed(inSpriteXValue_23) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_722 = {{1{inSpriteXValue_23[11]}},inSpriteXValue_23}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_940 = {{1{spriteYPositionReg_23[9]}},spriteYPositionReg_23}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_23 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_940); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_23 = inSpriteYValue_23[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_23 = $signed(inSpriteYPreScaled_23) >= 11'sh0 & $signed(inSpriteYPreScaled_23) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_730 = {{1{inSpriteYPreScaled_23[10]}},inSpriteYPreScaled_23}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_24 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_24); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_24 = $signed(inSpriteXValue_24) >= 12'sh0 & $signed(inSpriteXValue_24) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_738 = {{1{inSpriteXValue_24[11]}},inSpriteXValue_24}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_942 = {{1{spriteYPositionReg_24[9]}},spriteYPositionReg_24}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_24 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_942); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_24 = inSpriteYValue_24[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_24 = $signed(inSpriteYPreScaled_24) >= 11'sh0 & $signed(inSpriteYPreScaled_24) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_746 = {{1{inSpriteYPreScaled_24[10]}},inSpriteYPreScaled_24}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_25 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_25); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_25 = $signed(inSpriteXValue_25) >= 12'sh0 & $signed(inSpriteXValue_25) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_754 = {{1{inSpriteXValue_25[11]}},inSpriteXValue_25}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_944 = {{1{spriteYPositionReg_25[9]}},spriteYPositionReg_25}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_25 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_944); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_25 = inSpriteYValue_25[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_25 = $signed(inSpriteYPreScaled_25) >= 11'sh0 & $signed(inSpriteYPreScaled_25) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_762 = {{1{inSpriteYPreScaled_25[10]}},inSpriteYPreScaled_25}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_26 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_26); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_26 = $signed(inSpriteXValue_26) >= 12'sh0 & $signed(inSpriteXValue_26) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_770 = {{1{inSpriteXValue_26[11]}},inSpriteXValue_26}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_946 = {{1{spriteYPositionReg_26[9]}},spriteYPositionReg_26}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_26 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_946); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_26 = inSpriteYValue_26[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_26 = $signed(inSpriteYPreScaled_26) >= 11'sh0 & $signed(inSpriteYPreScaled_26) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_778 = {{1{inSpriteYPreScaled_26[10]}},inSpriteYPreScaled_26}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_27 = $signed(_inSpriteXValue_T_1) - $signed(spriteXPositionReg_27); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_27 = $signed(inSpriteXValue_27) >= 12'sh0 & $signed(inSpriteXValue_27) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_786 = {{1{inSpriteXValue_27[11]}},inSpriteXValue_27}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [10:0] _GEN_948 = {{1{spriteYPositionReg_27[9]}},spriteYPositionReg_27}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [11:0] inSpriteYValue_27 = $signed(_inSpriteYValue_T_1) - $signed(_GEN_948); // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_27 = inSpriteYValue_27[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_27 = $signed(inSpriteYPreScaled_27) >= 11'sh0 & $signed(inSpriteYPreScaled_27) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_794 = {{1{inSpriteYPreScaled_27[10]}},inSpriteYPreScaled_27}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteXValue_28 = $signed(_inSpriteXValue_T_1) - 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 263:54]
  wire  inSpriteHorizontal_28 = $signed(inSpriteXValue_28) >= 12'sh0 & $signed(inSpriteXValue_28) < 12'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 272:61]
  wire [12:0] _GEN_802 = {{1{inSpriteXValue_28[11]}},inSpriteXValue_28}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 269:149 271:20]
  wire [11:0] inSpriteYValue_28 = $signed(_inSpriteYValue_T_1) - 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 292:54]
  wire [10:0] inSpriteYPreScaled_28 = inSpriteYValue_28[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 258:32]
  wire  inSpriteVertical_28 = $signed(inSpriteYPreScaled_28) >= 11'sh0 & $signed(inSpriteYPreScaled_28) < 11'sh20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 301:59]
  wire [11:0] _GEN_810 = {{1{inSpriteYPreScaled_28[10]}},inSpriteYPreScaled_28}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 298:142 300:20]
  wire [11:0] inSpriteX_0 = _GEN_354[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_0 = _GEN_362[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_0_io_address_T_2 = 6'h20 * inSpriteY_0[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_956 = {{6'd0}, inSpriteX_0[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_0_io_address_T_4 = _GEN_956 + _spriteMemories_0_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_1 = _GEN_370[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_1 = _GEN_378[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_1_io_address_T_2 = 6'h20 * inSpriteY_1[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_959 = {{6'd0}, inSpriteX_1[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_1_io_address_T_4 = _GEN_959 + _spriteMemories_1_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_2 = _GEN_386[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_2 = _GEN_394[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_2_io_address_T_2 = 6'h20 * inSpriteY_2[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_962 = {{6'd0}, inSpriteX_2[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_2_io_address_T_4 = _GEN_962 + _spriteMemories_2_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_3 = _GEN_402[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_3 = _GEN_410[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_3_io_address_T_2 = 6'h20 * inSpriteY_3[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_965 = {{6'd0}, inSpriteX_3[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_3_io_address_T_4 = _GEN_965 + _spriteMemories_3_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_4 = _GEN_418[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_4 = _GEN_426[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_4_io_address_T_2 = 6'h20 * inSpriteY_4[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_968 = {{6'd0}, inSpriteX_4[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_4_io_address_T_4 = _GEN_968 + _spriteMemories_4_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_5 = _GEN_434[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_5 = _GEN_442[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_5_io_address_T_2 = 6'h20 * inSpriteY_5[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_971 = {{6'd0}, inSpriteX_5[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_5_io_address_T_4 = _GEN_971 + _spriteMemories_5_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_6 = _GEN_450[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_6 = _GEN_458[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_6_io_address_T_2 = 6'h20 * inSpriteY_6[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_974 = {{6'd0}, inSpriteX_6[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_6_io_address_T_4 = _GEN_974 + _spriteMemories_6_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_7 = _GEN_466[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_7 = _GEN_474[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_7_io_address_T_2 = 6'h20 * inSpriteY_7[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_977 = {{6'd0}, inSpriteX_7[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_7_io_address_T_4 = _GEN_977 + _spriteMemories_7_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_8 = _GEN_482[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_8 = _GEN_490[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_8_io_address_T_2 = 6'h20 * inSpriteY_8[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_980 = {{6'd0}, inSpriteX_8[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_8_io_address_T_4 = _GEN_980 + _spriteMemories_8_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_9 = _GEN_498[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_9 = _GEN_506[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_9_io_address_T_2 = 6'h20 * inSpriteY_9[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_983 = {{6'd0}, inSpriteX_9[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_9_io_address_T_4 = _GEN_983 + _spriteMemories_9_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_10 = _GEN_514[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_10 = _GEN_522[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_10_io_address_T_2 = 6'h20 * inSpriteY_10[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_986 = {{6'd0}, inSpriteX_10[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_10_io_address_T_4 = _GEN_986 + _spriteMemories_10_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_11 = _GEN_530[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_11 = _GEN_538[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_11_io_address_T_2 = 6'h20 * inSpriteY_11[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_989 = {{6'd0}, inSpriteX_11[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_11_io_address_T_4 = _GEN_989 + _spriteMemories_11_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_12 = _GEN_546[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_12 = _GEN_554[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_12_io_address_T_2 = 6'h20 * inSpriteY_12[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_992 = {{6'd0}, inSpriteX_12[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_12_io_address_T_4 = _GEN_992 + _spriteMemories_12_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_13 = _GEN_562[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_13 = _GEN_570[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_13_io_address_T_2 = 6'h20 * inSpriteY_13[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_995 = {{6'd0}, inSpriteX_13[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_13_io_address_T_4 = _GEN_995 + _spriteMemories_13_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_14 = _GEN_578[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_14 = _GEN_586[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_14_io_address_T_2 = 6'h20 * inSpriteY_14[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_998 = {{6'd0}, inSpriteX_14[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_14_io_address_T_4 = _GEN_998 + _spriteMemories_14_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_15 = _GEN_594[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_15 = _GEN_602[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_15_io_address_T_2 = 6'h20 * inSpriteY_15[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1001 = {{6'd0}, inSpriteX_15[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_15_io_address_T_4 = _GEN_1001 + _spriteMemories_15_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_16 = _GEN_610[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_16 = _GEN_618[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_16_io_address_T_2 = 6'h20 * inSpriteY_16[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1004 = {{6'd0}, inSpriteX_16[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_16_io_address_T_4 = _GEN_1004 + _spriteMemories_16_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_17 = _GEN_626[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_17 = _GEN_634[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_17_io_address_T_2 = 6'h20 * inSpriteY_17[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1007 = {{6'd0}, inSpriteX_17[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_17_io_address_T_4 = _GEN_1007 + _spriteMemories_17_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_18 = _GEN_642[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_18 = _GEN_650[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_18_io_address_T_2 = 6'h20 * inSpriteY_18[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1010 = {{6'd0}, inSpriteX_18[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_18_io_address_T_4 = _GEN_1010 + _spriteMemories_18_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_19 = _GEN_658[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_19 = _GEN_666[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_19_io_address_T_2 = 6'h20 * inSpriteY_19[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1013 = {{6'd0}, inSpriteX_19[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_19_io_address_T_4 = _GEN_1013 + _spriteMemories_19_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_20 = _GEN_674[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_20 = _GEN_682[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_20_io_address_T_2 = 6'h20 * inSpriteY_20[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1016 = {{6'd0}, inSpriteX_20[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_20_io_address_T_4 = _GEN_1016 + _spriteMemories_20_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_21 = _GEN_690[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_21 = _GEN_698[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_21_io_address_T_2 = 6'h20 * inSpriteY_21[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1019 = {{6'd0}, inSpriteX_21[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_21_io_address_T_4 = _GEN_1019 + _spriteMemories_21_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_22 = _GEN_706[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_22 = _GEN_714[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_22_io_address_T_2 = 6'h20 * inSpriteY_22[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1022 = {{6'd0}, inSpriteX_22[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_22_io_address_T_4 = _GEN_1022 + _spriteMemories_22_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_23 = _GEN_722[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_23 = _GEN_730[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_23_io_address_T_2 = 6'h20 * inSpriteY_23[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1025 = {{6'd0}, inSpriteX_23[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_23_io_address_T_4 = _GEN_1025 + _spriteMemories_23_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_24 = _GEN_738[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_24 = _GEN_746[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_24_io_address_T_2 = 6'h20 * inSpriteY_24[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1028 = {{6'd0}, inSpriteX_24[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_24_io_address_T_4 = _GEN_1028 + _spriteMemories_24_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_25 = _GEN_754[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_25 = _GEN_762[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_25_io_address_T_2 = 6'h20 * inSpriteY_25[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1031 = {{6'd0}, inSpriteX_25[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_25_io_address_T_4 = _GEN_1031 + _spriteMemories_25_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_26 = _GEN_770[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_26 = _GEN_778[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_26_io_address_T_2 = 6'h20 * inSpriteY_26[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1034 = {{6'd0}, inSpriteX_26[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_26_io_address_T_4 = _GEN_1034 + _spriteMemories_26_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_27 = _GEN_786[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_27 = _GEN_794[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_27_io_address_T_2 = 6'h20 * inSpriteY_27[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1037 = {{6'd0}, inSpriteX_27[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_27_io_address_T_4 = _GEN_1037 + _spriteMemories_27_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [11:0] inSpriteX_28 = _GEN_802[11:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 259:23]
  wire [10:0] inSpriteY_28 = _GEN_810[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 260:23]
  wire [10:0] _spriteMemories_28_io_address_T_2 = 6'h20 * inSpriteY_28[4:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:74]
  wire [10:0] _GEN_1040 = {{6'd0}, inSpriteX_28[4:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  wire [10:0] _spriteMemories_28_io_address_T_4 = _GEN_1040 + _spriteMemories_28_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:62]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] multiHotPriortyReductionTree_io_dataInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:60]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  multiHotPriortyReductionTree_io_selectInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:132]
  reg [5:0] pixelColorSprite; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 339:33]
  reg  pixelColorSpriteValid; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 340:38]
  wire [5:0] pixelColorInDisplay = pixelColorSpriteValid ? pixelColorSprite : pixelColorBack; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 344:32]
  reg  pixelColourVGA_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  pixelColourVGA_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  reg  pixelColourVGA_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 21:24]
  wire [5:0] pixelColourVGA = pixelColourVGA_pipeReg_0 ? pixelColorInDisplay : 6'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 345:27]
  reg [3:0] io_vgaRed_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 349:23]
  reg [3:0] io_vgaGreen_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 350:25]
  reg [3:0] io_vgaBlue_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 351:24]
  Memory backTileMemories_0 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_0_clock),
    .io_address(backTileMemories_0_io_address),
    .io_dataRead(backTileMemories_0_io_dataRead)
  );
  Memory_1 backTileMemories_1 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_1_clock),
    .io_address(backTileMemories_1_io_address),
    .io_dataRead(backTileMemories_1_io_dataRead)
  );
  Memory_2 backTileMemories_2 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_2_clock),
    .io_address(backTileMemories_2_io_address),
    .io_dataRead(backTileMemories_2_io_dataRead)
  );
  Memory_3 backTileMemories_3 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_3_clock),
    .io_address(backTileMemories_3_io_address),
    .io_dataRead(backTileMemories_3_io_dataRead)
  );
  Memory_4 backTileMemories_4 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_4_clock),
    .io_address(backTileMemories_4_io_address),
    .io_dataRead(backTileMemories_4_io_dataRead)
  );
  Memory_5 backTileMemories_5 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_5_clock),
    .io_address(backTileMemories_5_io_address),
    .io_dataRead(backTileMemories_5_io_dataRead)
  );
  Memory_6 backTileMemories_6 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_6_clock),
    .io_address(backTileMemories_6_io_address),
    .io_dataRead(backTileMemories_6_io_dataRead)
  );
  Memory_7 backTileMemories_7 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_7_clock),
    .io_address(backTileMemories_7_io_address),
    .io_dataRead(backTileMemories_7_io_dataRead)
  );
  Memory_8 backTileMemories_8 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_8_clock),
    .io_address(backTileMemories_8_io_address),
    .io_dataRead(backTileMemories_8_io_dataRead)
  );
  Memory_9 backTileMemories_9 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_9_clock),
    .io_address(backTileMemories_9_io_address),
    .io_dataRead(backTileMemories_9_io_dataRead)
  );
  Memory_10 backTileMemories_10 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_10_clock),
    .io_address(backTileMemories_10_io_address),
    .io_dataRead(backTileMemories_10_io_dataRead)
  );
  Memory_11 backTileMemories_11 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_11_clock),
    .io_address(backTileMemories_11_io_address),
    .io_dataRead(backTileMemories_11_io_dataRead)
  );
  Memory_12 backTileMemories_12 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_12_clock),
    .io_address(backTileMemories_12_io_address),
    .io_dataRead(backTileMemories_12_io_dataRead)
  );
  Memory_13 backTileMemories_13 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_13_clock),
    .io_address(backTileMemories_13_io_address),
    .io_dataRead(backTileMemories_13_io_dataRead)
  );
  Memory_14 backTileMemories_14 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_14_clock),
    .io_address(backTileMemories_14_io_address),
    .io_dataRead(backTileMemories_14_io_dataRead)
  );
  Memory_15 backTileMemories_15 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_15_clock),
    .io_address(backTileMemories_15_io_address),
    .io_dataRead(backTileMemories_15_io_dataRead)
  );
  Memory_16 backTileMemories_16 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_16_clock),
    .io_address(backTileMemories_16_io_address),
    .io_dataRead(backTileMemories_16_io_dataRead)
  );
  Memory_17 backTileMemories_17 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_17_clock),
    .io_address(backTileMemories_17_io_address),
    .io_dataRead(backTileMemories_17_io_dataRead)
  );
  Memory_18 backTileMemories_18 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_18_clock),
    .io_address(backTileMemories_18_io_address),
    .io_dataRead(backTileMemories_18_io_dataRead)
  );
  Memory_19 backTileMemories_19 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_19_clock),
    .io_address(backTileMemories_19_io_address),
    .io_dataRead(backTileMemories_19_io_dataRead)
  );
  Memory_20 backTileMemories_20 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_20_clock),
    .io_address(backTileMemories_20_io_address),
    .io_dataRead(backTileMemories_20_io_dataRead)
  );
  Memory_21 backTileMemories_21 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_21_clock),
    .io_address(backTileMemories_21_io_address),
    .io_dataRead(backTileMemories_21_io_dataRead)
  );
  Memory_22 backTileMemories_22 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_22_clock),
    .io_address(backTileMemories_22_io_address),
    .io_dataRead(backTileMemories_22_io_dataRead)
  );
  Memory_23 backTileMemories_23 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_23_clock),
    .io_address(backTileMemories_23_io_address),
    .io_dataRead(backTileMemories_23_io_dataRead)
  );
  Memory_24 backTileMemories_24 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_24_clock),
    .io_address(backTileMemories_24_io_address),
    .io_dataRead(backTileMemories_24_io_dataRead)
  );
  Memory_25 backTileMemories_25 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_25_clock),
    .io_address(backTileMemories_25_io_address),
    .io_dataRead(backTileMemories_25_io_dataRead)
  );
  Memory_26 backTileMemories_26 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_26_clock),
    .io_address(backTileMemories_26_io_address),
    .io_dataRead(backTileMemories_26_io_dataRead)
  );
  Memory_27 backTileMemories_27 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_27_clock),
    .io_address(backTileMemories_27_io_address),
    .io_dataRead(backTileMemories_27_io_dataRead)
  );
  Memory_28 backTileMemories_28 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_28_clock),
    .io_address(backTileMemories_28_io_address),
    .io_dataRead(backTileMemories_28_io_dataRead)
  );
  Memory_29 backTileMemories_29 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_29_clock),
    .io_address(backTileMemories_29_io_address),
    .io_dataRead(backTileMemories_29_io_dataRead)
  );
  Memory_30 backTileMemories_30 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_30_clock),
    .io_address(backTileMemories_30_io_address),
    .io_dataRead(backTileMemories_30_io_dataRead)
  );
  Memory_31 backTileMemories_31 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 161:32]
    .clock(backTileMemories_31_clock),
    .io_address(backTileMemories_31_io_address),
    .io_dataRead(backTileMemories_31_io_dataRead)
  );
  Memory_32 backBufferMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 178:32]
    .clock(backBufferMemory_clock),
    .io_address(backBufferMemory_io_address),
    .io_dataRead(backBufferMemory_io_dataRead),
    .io_writeEnable(backBufferMemory_io_writeEnable),
    .io_dataWrite(backBufferMemory_io_dataWrite)
  );
  Memory_32 backBufferShadowMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 179:38]
    .clock(backBufferShadowMemory_clock),
    .io_address(backBufferShadowMemory_io_address),
    .io_dataRead(backBufferShadowMemory_io_dataRead),
    .io_writeEnable(backBufferShadowMemory_io_writeEnable),
    .io_dataWrite(backBufferShadowMemory_io_dataWrite)
  );
  Memory_34 backBufferRestoreMemory ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 180:39]
    .clock(backBufferRestoreMemory_clock),
    .io_address(backBufferRestoreMemory_io_address),
    .io_dataRead(backBufferRestoreMemory_io_dataRead)
  );
  Memory_35 spriteMemories_0 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_0_clock),
    .io_address(spriteMemories_0_io_address),
    .io_dataRead(spriteMemories_0_io_dataRead)
  );
  Memory_36 spriteMemories_1 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_1_clock),
    .io_address(spriteMemories_1_io_address),
    .io_dataRead(spriteMemories_1_io_dataRead)
  );
  Memory_37 spriteMemories_2 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_2_clock),
    .io_address(spriteMemories_2_io_address),
    .io_dataRead(spriteMemories_2_io_dataRead)
  );
  Memory_38 spriteMemories_3 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_3_clock),
    .io_address(spriteMemories_3_io_address),
    .io_dataRead(spriteMemories_3_io_dataRead)
  );
  Memory_39 spriteMemories_4 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_4_clock),
    .io_address(spriteMemories_4_io_address),
    .io_dataRead(spriteMemories_4_io_dataRead)
  );
  Memory_40 spriteMemories_5 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_5_clock),
    .io_address(spriteMemories_5_io_address),
    .io_dataRead(spriteMemories_5_io_dataRead)
  );
  Memory_41 spriteMemories_6 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_6_clock),
    .io_address(spriteMemories_6_io_address),
    .io_dataRead(spriteMemories_6_io_dataRead)
  );
  Memory_42 spriteMemories_7 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_7_clock),
    .io_address(spriteMemories_7_io_address),
    .io_dataRead(spriteMemories_7_io_dataRead)
  );
  Memory_43 spriteMemories_8 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_8_clock),
    .io_address(spriteMemories_8_io_address),
    .io_dataRead(spriteMemories_8_io_dataRead)
  );
  Memory_44 spriteMemories_9 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_9_clock),
    .io_address(spriteMemories_9_io_address),
    .io_dataRead(spriteMemories_9_io_dataRead)
  );
  Memory_45 spriteMemories_10 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_10_clock),
    .io_address(spriteMemories_10_io_address),
    .io_dataRead(spriteMemories_10_io_dataRead)
  );
  Memory_46 spriteMemories_11 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_11_clock),
    .io_address(spriteMemories_11_io_address),
    .io_dataRead(spriteMemories_11_io_dataRead)
  );
  Memory_47 spriteMemories_12 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_12_clock),
    .io_address(spriteMemories_12_io_address),
    .io_dataRead(spriteMemories_12_io_dataRead)
  );
  Memory_48 spriteMemories_13 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_13_clock),
    .io_address(spriteMemories_13_io_address),
    .io_dataRead(spriteMemories_13_io_dataRead)
  );
  Memory_49 spriteMemories_14 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_14_clock),
    .io_address(spriteMemories_14_io_address),
    .io_dataRead(spriteMemories_14_io_dataRead)
  );
  Memory_50 spriteMemories_15 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_15_clock),
    .io_address(spriteMemories_15_io_address),
    .io_dataRead(spriteMemories_15_io_dataRead)
  );
  Memory_51 spriteMemories_16 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_16_clock),
    .io_address(spriteMemories_16_io_address),
    .io_dataRead(spriteMemories_16_io_dataRead)
  );
  Memory_52 spriteMemories_17 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_17_clock),
    .io_address(spriteMemories_17_io_address),
    .io_dataRead(spriteMemories_17_io_dataRead)
  );
  Memory_53 spriteMemories_18 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_18_clock),
    .io_address(spriteMemories_18_io_address),
    .io_dataRead(spriteMemories_18_io_dataRead)
  );
  Memory_54 spriteMemories_19 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_19_clock),
    .io_address(spriteMemories_19_io_address),
    .io_dataRead(spriteMemories_19_io_dataRead)
  );
  Memory_55 spriteMemories_20 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_20_clock),
    .io_address(spriteMemories_20_io_address),
    .io_dataRead(spriteMemories_20_io_dataRead)
  );
  Memory_56 spriteMemories_21 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_21_clock),
    .io_address(spriteMemories_21_io_address),
    .io_dataRead(spriteMemories_21_io_dataRead)
  );
  Memory_57 spriteMemories_22 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_22_clock),
    .io_address(spriteMemories_22_io_address),
    .io_dataRead(spriteMemories_22_io_dataRead)
  );
  Memory_58 spriteMemories_23 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_23_clock),
    .io_address(spriteMemories_23_io_address),
    .io_dataRead(spriteMemories_23_io_dataRead)
  );
  Memory_59 spriteMemories_24 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_24_clock),
    .io_address(spriteMemories_24_io_address),
    .io_dataRead(spriteMemories_24_io_dataRead)
  );
  Memory_60 spriteMemories_25 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_25_clock),
    .io_address(spriteMemories_25_io_address),
    .io_dataRead(spriteMemories_25_io_dataRead)
  );
  Memory_61 spriteMemories_26 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_26_clock),
    .io_address(spriteMemories_26_io_address),
    .io_dataRead(spriteMemories_26_io_dataRead)
  );
  Memory_62 spriteMemories_27 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_27_clock),
    .io_address(spriteMemories_27_io_address),
    .io_dataRead(spriteMemories_27_io_dataRead)
  );
  Memory_63 spriteMemories_28 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_28_clock),
    .io_address(spriteMemories_28_io_address),
    .io_dataRead(spriteMemories_28_io_dataRead)
  );
  Memory_64 spriteMemories_29 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_29_clock),
    .io_address(spriteMemories_29_io_address),
    .io_dataRead(spriteMemories_29_io_dataRead)
  );
  Memory_65 spriteMemories_30 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_30_clock),
    .io_address(spriteMemories_30_io_address),
    .io_dataRead(spriteMemories_30_io_dataRead)
  );
  Memory_66 spriteMemories_31 ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 250:30]
    .clock(spriteMemories_31_clock),
    .io_address(spriteMemories_31_io_address),
    .io_dataRead(spriteMemories_31_io_dataRead)
  );
  MultiHotPriortyReductionTree multiHotPriortyReductionTree ( // @[\\src\\main\\scala\\GraphicEngineVGA.scala 334:44]
    .io_dataInput_0(multiHotPriortyReductionTree_io_dataInput_0),
    .io_dataInput_1(multiHotPriortyReductionTree_io_dataInput_1),
    .io_dataInput_2(multiHotPriortyReductionTree_io_dataInput_2),
    .io_dataInput_3(multiHotPriortyReductionTree_io_dataInput_3),
    .io_dataInput_4(multiHotPriortyReductionTree_io_dataInput_4),
    .io_dataInput_5(multiHotPriortyReductionTree_io_dataInput_5),
    .io_dataInput_6(multiHotPriortyReductionTree_io_dataInput_6),
    .io_dataInput_7(multiHotPriortyReductionTree_io_dataInput_7),
    .io_dataInput_8(multiHotPriortyReductionTree_io_dataInput_8),
    .io_dataInput_9(multiHotPriortyReductionTree_io_dataInput_9),
    .io_dataInput_10(multiHotPriortyReductionTree_io_dataInput_10),
    .io_dataInput_11(multiHotPriortyReductionTree_io_dataInput_11),
    .io_dataInput_12(multiHotPriortyReductionTree_io_dataInput_12),
    .io_dataInput_13(multiHotPriortyReductionTree_io_dataInput_13),
    .io_dataInput_14(multiHotPriortyReductionTree_io_dataInput_14),
    .io_dataInput_15(multiHotPriortyReductionTree_io_dataInput_15),
    .io_dataInput_16(multiHotPriortyReductionTree_io_dataInput_16),
    .io_dataInput_17(multiHotPriortyReductionTree_io_dataInput_17),
    .io_dataInput_18(multiHotPriortyReductionTree_io_dataInput_18),
    .io_dataInput_19(multiHotPriortyReductionTree_io_dataInput_19),
    .io_dataInput_20(multiHotPriortyReductionTree_io_dataInput_20),
    .io_dataInput_21(multiHotPriortyReductionTree_io_dataInput_21),
    .io_dataInput_22(multiHotPriortyReductionTree_io_dataInput_22),
    .io_dataInput_23(multiHotPriortyReductionTree_io_dataInput_23),
    .io_dataInput_24(multiHotPriortyReductionTree_io_dataInput_24),
    .io_dataInput_25(multiHotPriortyReductionTree_io_dataInput_25),
    .io_dataInput_26(multiHotPriortyReductionTree_io_dataInput_26),
    .io_dataInput_27(multiHotPriortyReductionTree_io_dataInput_27),
    .io_dataInput_28(multiHotPriortyReductionTree_io_dataInput_28),
    .io_dataInput_29(multiHotPriortyReductionTree_io_dataInput_29),
    .io_dataInput_30(multiHotPriortyReductionTree_io_dataInput_30),
    .io_dataInput_31(multiHotPriortyReductionTree_io_dataInput_31),
    .io_selectInput_0(multiHotPriortyReductionTree_io_selectInput_0),
    .io_selectInput_1(multiHotPriortyReductionTree_io_selectInput_1),
    .io_selectInput_2(multiHotPriortyReductionTree_io_selectInput_2),
    .io_selectInput_3(multiHotPriortyReductionTree_io_selectInput_3),
    .io_selectInput_4(multiHotPriortyReductionTree_io_selectInput_4),
    .io_selectInput_5(multiHotPriortyReductionTree_io_selectInput_5),
    .io_selectInput_6(multiHotPriortyReductionTree_io_selectInput_6),
    .io_selectInput_7(multiHotPriortyReductionTree_io_selectInput_7),
    .io_selectInput_8(multiHotPriortyReductionTree_io_selectInput_8),
    .io_selectInput_9(multiHotPriortyReductionTree_io_selectInput_9),
    .io_selectInput_10(multiHotPriortyReductionTree_io_selectInput_10),
    .io_selectInput_11(multiHotPriortyReductionTree_io_selectInput_11),
    .io_selectInput_12(multiHotPriortyReductionTree_io_selectInput_12),
    .io_selectInput_13(multiHotPriortyReductionTree_io_selectInput_13),
    .io_selectInput_14(multiHotPriortyReductionTree_io_selectInput_14),
    .io_selectInput_15(multiHotPriortyReductionTree_io_selectInput_15),
    .io_selectInput_16(multiHotPriortyReductionTree_io_selectInput_16),
    .io_selectInput_17(multiHotPriortyReductionTree_io_selectInput_17),
    .io_selectInput_18(multiHotPriortyReductionTree_io_selectInput_18),
    .io_selectInput_19(multiHotPriortyReductionTree_io_selectInput_19),
    .io_selectInput_20(multiHotPriortyReductionTree_io_selectInput_20),
    .io_selectInput_21(multiHotPriortyReductionTree_io_selectInput_21),
    .io_selectInput_22(multiHotPriortyReductionTree_io_selectInput_22),
    .io_selectInput_23(multiHotPriortyReductionTree_io_selectInput_23),
    .io_selectInput_24(multiHotPriortyReductionTree_io_selectInput_24),
    .io_selectInput_25(multiHotPriortyReductionTree_io_selectInput_25),
    .io_selectInput_26(multiHotPriortyReductionTree_io_selectInput_26),
    .io_selectInput_27(multiHotPriortyReductionTree_io_selectInput_27),
    .io_selectInput_28(multiHotPriortyReductionTree_io_selectInput_28),
    .io_selectInput_29(multiHotPriortyReductionTree_io_selectInput_29),
    .io_selectInput_30(multiHotPriortyReductionTree_io_selectInput_30),
    .io_selectInput_31(multiHotPriortyReductionTree_io_selectInput_31),
    .io_dataOutput(multiHotPriortyReductionTree_io_dataOutput),
    .io_selectOutput(multiHotPriortyReductionTree_io_selectOutput)
  );
  assign io_newFrame = run & _GEN_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13 71:15]
  assign io_missingFrameError = missingFrameErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 131:24]
  assign io_backBufferWriteError = backBufferWriteErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 132:27]
  assign io_viewBoxOutOfRangeError = viewBoxOutOfRangeErrorReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 133:29]
  assign io_vgaRed = io_vgaRed_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 349:13]
  assign io_vgaBlue = io_vgaBlue_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 351:14]
  assign io_vgaGreen = io_vgaGreen_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 350:15]
  assign io_Hsync = io_Hsync_pipeReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 94:12]
  assign io_Vsync = io_Vsync_pipeReg_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 95:12]
  assign backTileMemories_0_clock = clock;
  assign backTileMemories_0_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_1_clock = clock;
  assign backTileMemories_1_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_2_clock = clock;
  assign backTileMemories_2_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_3_clock = clock;
  assign backTileMemories_3_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_4_clock = clock;
  assign backTileMemories_4_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_5_clock = clock;
  assign backTileMemories_5_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_6_clock = clock;
  assign backTileMemories_6_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_7_clock = clock;
  assign backTileMemories_7_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_8_clock = clock;
  assign backTileMemories_8_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_9_clock = clock;
  assign backTileMemories_9_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_10_clock = clock;
  assign backTileMemories_10_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_11_clock = clock;
  assign backTileMemories_11_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_12_clock = clock;
  assign backTileMemories_12_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_13_clock = clock;
  assign backTileMemories_13_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_14_clock = clock;
  assign backTileMemories_14_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_15_clock = clock;
  assign backTileMemories_15_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_16_clock = clock;
  assign backTileMemories_16_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_17_clock = clock;
  assign backTileMemories_17_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_18_clock = clock;
  assign backTileMemories_18_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_19_clock = clock;
  assign backTileMemories_19_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_20_clock = clock;
  assign backTileMemories_20_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_21_clock = clock;
  assign backTileMemories_21_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_22_clock = clock;
  assign backTileMemories_22_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_23_clock = clock;
  assign backTileMemories_23_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_24_clock = clock;
  assign backTileMemories_24_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_25_clock = clock;
  assign backTileMemories_25_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_26_clock = clock;
  assign backTileMemories_26_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_27_clock = clock;
  assign backTileMemories_27_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_28_clock = clock;
  assign backTileMemories_28_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_29_clock = clock;
  assign backTileMemories_29_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_30_clock = clock;
  assign backTileMemories_30_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backTileMemories_31_clock = clock;
  assign backTileMemories_31_io_address = _backTileMemories_0_io_address_T_3[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 172:36]
  assign backBufferMemory_clock = clock;
  assign backBufferMemory_io_address = _backBufferMemory_io_address_T_5[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:31]
  assign backBufferMemory_io_writeEnable = copyEnabledReg; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 228:35]
  assign backBufferMemory_io_dataWrite = backBufferShadowMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 229:33]
  assign backBufferShadowMemory_clock = clock;
  assign backBufferShadowMemory_io_address = restoreEnabled ? backBufferShadowMemory_io_address_REG :
    _backBufferShadowMemory_io_address_T_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:43]
  assign backBufferShadowMemory_io_writeEnable = restoreEnabled ? backBufferShadowMemory_io_writeEnable_REG :
    _backBufferShadowMemory_io_writeEnable_T; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:47]
  assign backBufferShadowMemory_io_dataWrite = restoreEnabled ? backBufferRestoreMemory_io_dataRead :
    backBufferShadowMemory_io_dataWrite_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 224:45]
  assign backBufferRestoreMemory_clock = clock;
  assign backBufferRestoreMemory_io_address = backMemoryRestoreCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 216:65]
  assign spriteMemories_0_clock = clock;
  assign spriteMemories_0_io_address = _spriteMemories_0_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_1_clock = clock;
  assign spriteMemories_1_io_address = _spriteMemories_1_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_2_clock = clock;
  assign spriteMemories_2_io_address = _spriteMemories_2_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_3_clock = clock;
  assign spriteMemories_3_io_address = _spriteMemories_3_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_4_clock = clock;
  assign spriteMemories_4_io_address = _spriteMemories_4_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_5_clock = clock;
  assign spriteMemories_5_io_address = _spriteMemories_5_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_6_clock = clock;
  assign spriteMemories_6_io_address = _spriteMemories_6_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_7_clock = clock;
  assign spriteMemories_7_io_address = _spriteMemories_7_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_8_clock = clock;
  assign spriteMemories_8_io_address = _spriteMemories_8_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_9_clock = clock;
  assign spriteMemories_9_io_address = _spriteMemories_9_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_10_clock = clock;
  assign spriteMemories_10_io_address = _spriteMemories_10_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_11_clock = clock;
  assign spriteMemories_11_io_address = _spriteMemories_11_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_12_clock = clock;
  assign spriteMemories_12_io_address = _spriteMemories_12_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_13_clock = clock;
  assign spriteMemories_13_io_address = _spriteMemories_13_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_14_clock = clock;
  assign spriteMemories_14_io_address = _spriteMemories_14_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_15_clock = clock;
  assign spriteMemories_15_io_address = _spriteMemories_15_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_16_clock = clock;
  assign spriteMemories_16_io_address = _spriteMemories_16_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_17_clock = clock;
  assign spriteMemories_17_io_address = _spriteMemories_17_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_18_clock = clock;
  assign spriteMemories_18_io_address = _spriteMemories_18_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_19_clock = clock;
  assign spriteMemories_19_io_address = _spriteMemories_19_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_20_clock = clock;
  assign spriteMemories_20_io_address = _spriteMemories_20_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_21_clock = clock;
  assign spriteMemories_21_io_address = _spriteMemories_21_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_22_clock = clock;
  assign spriteMemories_22_io_address = _spriteMemories_22_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_23_clock = clock;
  assign spriteMemories_23_io_address = _spriteMemories_23_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_24_clock = clock;
  assign spriteMemories_24_io_address = _spriteMemories_24_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_25_clock = clock;
  assign spriteMemories_25_io_address = _spriteMemories_25_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_26_clock = clock;
  assign spriteMemories_26_io_address = _spriteMemories_26_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_27_clock = clock;
  assign spriteMemories_27_io_address = _spriteMemories_27_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_28_clock = clock;
  assign spriteMemories_28_io_address = _spriteMemories_28_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_29_clock = clock;
  assign spriteMemories_29_io_address = _spriteMemories_28_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_30_clock = clock;
  assign spriteMemories_30_io_address = _spriteMemories_28_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign spriteMemories_31_clock = clock;
  assign spriteMemories_31_io_address = _spriteMemories_28_io_address_T_4[9:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 329:34]
  assign multiHotPriortyReductionTree_io_dataInput_0 = multiHotPriortyReductionTree_io_dataInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_1 = multiHotPriortyReductionTree_io_dataInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_2 = multiHotPriortyReductionTree_io_dataInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_3 = multiHotPriortyReductionTree_io_dataInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_4 = multiHotPriortyReductionTree_io_dataInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_5 = multiHotPriortyReductionTree_io_dataInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_6 = multiHotPriortyReductionTree_io_dataInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_7 = multiHotPriortyReductionTree_io_dataInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_8 = multiHotPriortyReductionTree_io_dataInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_9 = multiHotPriortyReductionTree_io_dataInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_10 = multiHotPriortyReductionTree_io_dataInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_11 = multiHotPriortyReductionTree_io_dataInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_12 = multiHotPriortyReductionTree_io_dataInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_13 = multiHotPriortyReductionTree_io_dataInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_14 = multiHotPriortyReductionTree_io_dataInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_15 = multiHotPriortyReductionTree_io_dataInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_16 = multiHotPriortyReductionTree_io_dataInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_17 = multiHotPriortyReductionTree_io_dataInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_18 = multiHotPriortyReductionTree_io_dataInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_19 = multiHotPriortyReductionTree_io_dataInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_20 = multiHotPriortyReductionTree_io_dataInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_21 = multiHotPriortyReductionTree_io_dataInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_22 = multiHotPriortyReductionTree_io_dataInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_23 = multiHotPriortyReductionTree_io_dataInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_24 = multiHotPriortyReductionTree_io_dataInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_25 = multiHotPriortyReductionTree_io_dataInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_26 = multiHotPriortyReductionTree_io_dataInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_27 = multiHotPriortyReductionTree_io_dataInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_28 = multiHotPriortyReductionTree_io_dataInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_29 = multiHotPriortyReductionTree_io_dataInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_30 = multiHotPriortyReductionTree_io_dataInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_dataInput_31 = multiHotPriortyReductionTree_io_dataInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:50]
  assign multiHotPriortyReductionTree_io_selectInput_0 = multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_0_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_1 = multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_1_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_2 = multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_2_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_3 = multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_3_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_4 = multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_4_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_5 = multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_5_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_6 = multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_6_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_7 = multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_7_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_8 = multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_8_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_9 = multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_9_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_10 = multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_10_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_11 = multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_11_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_12 = multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_12_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_13 = multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_13_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_14 = multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_14_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_15 = multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_15_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_16 = multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_16_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_17 = multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_17_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_18 = multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_18_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_19 = multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_19_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_20 = multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_20_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_21 = multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_21_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_22 = multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_22_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_23 = multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_23_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_24 = multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_24_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_25 = multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_25_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_26 = multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_26_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_27 = multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_27_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_28 = multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_28_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_29 = multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_29_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_30 = multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_30_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  assign multiHotPriortyReductionTree_io_selectInput_31 = multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 &
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 & ~multiHotPriortyReductionTree_io_selectInput_31_REG; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:121]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
      ScaleCounterReg <= 2'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 67:32]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        ScaleCounterReg <= 2'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 75:23]
      end else begin
        ScaleCounterReg <= _ScaleCounterReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 88:23]
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
      CounterXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 68:28]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        if (CounterXReg == 10'h31f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129]
          CounterXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 77:21]
        end else begin
          CounterXReg <= _CounterXReg_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 85:21]
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
      CounterYReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 69:28]
    end else if (run) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 73:13]
      if (ScaleCounterReg == 2'h3) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 74:52]
        if (CounterXReg == 10'h31f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 76:129]
          CounterYReg <= _GEN_0;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
      backMemoryRestoreCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 202:41]
    end else if (restoreEnabled) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:70]
      backMemoryRestoreCounter <= _backMemoryRestoreCounter_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 206:30]
    end
    io_Hsync_pipeReg_0 <= io_Hsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_1 <= io_Hsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_2 <= io_Hsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Hsync_pipeReg_3 <= ~Hsync; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 94:27]
    io_Vsync_pipeReg_0 <= io_Vsync_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_1 <= io_Vsync_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_2 <= io_Vsync_pipeReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    io_Vsync_pipeReg_3 <= ~Vsync; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 95:27]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
      frameClockCount <= 21'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 104:32]
    end else if (frameClockCount == 21'h19a27f) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 105:25]
      frameClockCount <= 21'h0;
    end else begin
      frameClockCount <= _frameClockCount_T_2;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_0 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_0 <= io_spriteXPosition_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_1 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_1 <= io_spriteXPosition_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_2 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_2 <= io_spriteXPosition_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_3 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_3 <= io_spriteXPosition_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_4 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_4 <= io_spriteXPosition_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_5 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_5 <= io_spriteXPosition_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_6 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_6 <= io_spriteXPosition_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_7 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_7 <= io_spriteXPosition_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_8 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_8 <= io_spriteXPosition_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_9 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_9 <= io_spriteXPosition_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_10 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_10 <= io_spriteXPosition_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_11 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_11 <= io_spriteXPosition_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_12 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_12 <= io_spriteXPosition_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_13 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_13 <= io_spriteXPosition_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_14 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_14 <= io_spriteXPosition_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_15 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_15 <= io_spriteXPosition_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_16 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_16 <= io_spriteXPosition_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_17 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_17 <= io_spriteXPosition_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_18 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_18 <= io_spriteXPosition_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_19 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_19 <= io_spriteXPosition_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_20 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_20 <= io_spriteXPosition_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_21 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_21 <= io_spriteXPosition_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_22 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_22 <= io_spriteXPosition_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_23 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_23 <= io_spriteXPosition_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_24 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_24 <= io_spriteXPosition_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_25 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_25 <= io_spriteXPosition_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_26 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_26 <= io_spriteXPosition_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_27 <= 11'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
      spriteXPositionReg_27 <= io_spriteXPosition_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 114:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_0 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_0 <= io_spriteYPosition_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_1 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_1 <= io_spriteYPosition_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_2 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_2 <= io_spriteYPosition_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_3 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_3 <= io_spriteYPosition_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_4 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_4 <= io_spriteYPosition_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_5 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_5 <= io_spriteYPosition_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_6 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_6 <= io_spriteYPosition_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_7 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_7 <= io_spriteYPosition_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_8 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_8 <= io_spriteYPosition_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_9 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_9 <= io_spriteYPosition_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_10 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_10 <= io_spriteYPosition_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_11 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_11 <= io_spriteYPosition_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_12 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_12 <= io_spriteYPosition_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_13 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_13 <= io_spriteYPosition_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_14 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_14 <= io_spriteYPosition_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_15 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_15 <= io_spriteYPosition_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_16 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_16 <= io_spriteYPosition_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_17 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_17 <= io_spriteYPosition_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_18 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_18 <= io_spriteYPosition_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_19 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_19 <= io_spriteYPosition_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_20 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_20 <= io_spriteYPosition_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_21 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_21 <= io_spriteYPosition_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_22 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_22 <= io_spriteYPosition_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_23 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_23 <= io_spriteYPosition_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_24 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_24 <= io_spriteYPosition_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_25 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_25 <= io_spriteYPosition_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_26 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_26 <= io_spriteYPosition_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_27 <= 10'sh0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
      spriteYPositionReg_27 <= io_spriteYPosition_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 115:37]
    end
    spriteVisibleReg_0 <= reset | _GEN_77; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_1 <= reset | _GEN_78; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_2 <= reset | _GEN_79; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_3 <= reset | _GEN_80; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_4 <= reset | _GEN_81; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_5 <= reset | _GEN_82; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_6 <= reset | _GEN_83; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_7 <= reset | _GEN_84; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_8 <= reset | _GEN_85; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_9 <= reset | _GEN_86; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_10 <= reset | _GEN_87; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_11 <= reset | _GEN_88; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_12 <= reset | _GEN_89; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_13 <= reset | _GEN_90; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_14 <= reset | _GEN_91; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_15 <= reset | _GEN_92; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_16 <= reset | _GEN_93; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_17 <= reset | _GEN_94; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_18 <= reset | _GEN_95; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_19 <= reset | _GEN_96; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_20 <= reset | _GEN_97; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_21 <= reset | _GEN_98; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_22 <= reset | _GEN_99; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_23 <= reset | _GEN_100; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_24 <= reset | _GEN_101; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_25 <= reset | _GEN_102; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_26 <= reset | _GEN_103; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_27 <= reset | _GEN_104; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_28 <= reset | _GEN_105; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_29 <= reset | _GEN_106; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_30 <= reset | _GEN_107; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    spriteVisibleReg_31 <= reset | _GEN_108; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 116:{35,35}]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
      viewBoxXReg <= io_viewBoxX; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 123:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
      viewBoxYReg <= 9'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
    end else if (io_newFrame) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
      viewBoxYReg <= io_viewBoxY; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 124:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
      missingFrameErrorReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 128:37]
    end else begin
      missingFrameErrorReg <= _GEN_306;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 129:40]
      backBufferWriteErrorReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 129:40]
    end else if (copyEnabled | copyEnabledReg) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 233:39]
      backBufferWriteErrorReg <= _GEN_314;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
      viewBoxOutOfRangeErrorReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 130:42]
    end else begin
      viewBoxOutOfRangeErrorReg <= _GEN_303;
    end
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
      newFrameStikyReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 147:33]
    end else if (REG) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:37]
      newFrameStikyReg <= 1'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 152:22]
    end else begin
      newFrameStikyReg <= _GEN_304;
    end
    REG <= io_frameUpdateDone; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 151:16]
    backTileMemoryDataRead_0_REG <= backTileMemories_0_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_1_REG <= backTileMemories_1_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_2_REG <= backTileMemories_2_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_3_REG <= backTileMemories_3_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_4_REG <= backTileMemories_4_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_5_REG <= backTileMemories_5_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_6_REG <= backTileMemories_6_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_7_REG <= backTileMemories_7_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_8_REG <= backTileMemories_8_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_9_REG <= backTileMemories_9_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_10_REG <= backTileMemories_10_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_11_REG <= backTileMemories_11_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_12_REG <= backTileMemories_12_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_13_REG <= backTileMemories_13_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_14_REG <= backTileMemories_14_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_15_REG <= backTileMemories_15_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_16_REG <= backTileMemories_16_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_17_REG <= backTileMemories_17_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_18_REG <= backTileMemories_18_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_19_REG <= backTileMemories_19_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_20_REG <= backTileMemories_20_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_21_REG <= backTileMemories_21_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_22_REG <= backTileMemories_22_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_23_REG <= backTileMemories_23_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_24_REG <= backTileMemories_24_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_25_REG <= backTileMemories_25_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_26_REG <= backTileMemories_26_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_27_REG <= backTileMemories_27_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_28_REG <= backTileMemories_28_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_29_REG <= backTileMemories_29_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_30_REG <= backTileMemories_30_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    backTileMemoryDataRead_31_REG <= backTileMemories_31_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 173:41]
    if (reset) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
      backMemoryCopyCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 183:38]
    end else if (preDisplayArea) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23]
      if (backMemoryCopyCounter < 12'h800) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 187:66]
        backMemoryCopyCounter <= _backMemoryCopyCounter_T_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 188:29]
      end
    end else begin
      backMemoryCopyCounter <= 12'h0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 197:27]
    end
    copyEnabledReg <= preDisplayArea & _T_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 186:23 198:17]
    backBufferShadowMemory_io_address_REG <= backMemoryRestoreCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:92]
    backBufferShadowMemory_io_address_REG_1 <= io_backBufferWriteAddress; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 221:156]
    backBufferShadowMemory_io_writeEnable_REG <= backMemoryRestoreCounter < 12'h800; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 205:33]
    backBufferShadowMemory_io_writeEnable_REG_1 <= io_backBufferWriteEnable; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 223:122]
    backBufferShadowMemory_io_dataWrite_REG <= io_backBufferWriteData; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 224:106]
    backBufferMemory_io_address_REG <= backMemoryCopyCounter[10:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 226:83]
    fullBackgroundColor_REG <= backBufferMemory_io_dataRead; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 243:56]
    if (fullBackgroundColor[6]) begin // @[\\src\\main\\scala\\GraphicEngineVGA.scala 244:25]
      pixelColorBack <= 6'h0;
    end else begin
      pixelColorBack <= fullBackgroundColor[5:0];
    end
    multiHotPriortyReductionTree_io_dataInput_0_REG <= spriteMemories_0_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1 <= spriteVisibleReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1 <= inSpriteHorizontal_0 & inSpriteVertical_0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_0_REG <= spriteMemories_0_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_1_REG <= spriteMemories_1_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1 <= spriteVisibleReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1 <= inSpriteHorizontal_1 & inSpriteVertical_1; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_1_REG <= spriteMemories_1_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_2_REG <= spriteMemories_2_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1 <= spriteVisibleReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1 <= inSpriteHorizontal_2 & inSpriteVertical_2; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_2_REG <= spriteMemories_2_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_3_REG <= spriteMemories_3_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1 <= spriteVisibleReg_3; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1 <= inSpriteHorizontal_3 & inSpriteVertical_3; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_3_REG <= spriteMemories_3_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_4_REG <= spriteMemories_4_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1 <= spriteVisibleReg_4; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1 <= inSpriteHorizontal_4 & inSpriteVertical_4; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_4_REG <= spriteMemories_4_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_5_REG <= spriteMemories_5_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1 <= spriteVisibleReg_5; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1 <= inSpriteHorizontal_5 & inSpriteVertical_5; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_5_REG <= spriteMemories_5_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_6_REG <= spriteMemories_6_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1 <= spriteVisibleReg_6; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1 <= inSpriteHorizontal_6 & inSpriteVertical_6; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_6_REG <= spriteMemories_6_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_7_REG <= spriteMemories_7_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1 <= spriteVisibleReg_7; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1 <= inSpriteHorizontal_7 & inSpriteVertical_7; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_7_REG <= spriteMemories_7_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_8_REG <= spriteMemories_8_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1 <= spriteVisibleReg_8; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1 <= inSpriteHorizontal_8 & inSpriteVertical_8; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_8_REG <= spriteMemories_8_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_9_REG <= spriteMemories_9_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 <= multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1
      ; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1 <= spriteVisibleReg_9; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1 <= inSpriteHorizontal_9 & inSpriteVertical_9; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_9_REG <= spriteMemories_9_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_10_REG <= spriteMemories_10_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1 <= spriteVisibleReg_10; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1 <= inSpriteHorizontal_10 & inSpriteVertical_10; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_10_REG <= spriteMemories_10_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_11_REG <= spriteMemories_11_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1 <= spriteVisibleReg_11; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1 <= inSpriteHorizontal_11 & inSpriteVertical_11; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_11_REG <= spriteMemories_11_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_12_REG <= spriteMemories_12_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1 <= spriteVisibleReg_12; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1 <= inSpriteHorizontal_12 & inSpriteVertical_12; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_12_REG <= spriteMemories_12_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_13_REG <= spriteMemories_13_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1 <= spriteVisibleReg_13; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1 <= inSpriteHorizontal_13 & inSpriteVertical_13; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_13_REG <= spriteMemories_13_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_14_REG <= spriteMemories_14_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1 <= spriteVisibleReg_14; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1 <= inSpriteHorizontal_14 & inSpriteVertical_14; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_14_REG <= spriteMemories_14_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_15_REG <= spriteMemories_15_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1 <= spriteVisibleReg_15; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1 <= inSpriteHorizontal_15 & inSpriteVertical_15; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_15_REG <= spriteMemories_15_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_16_REG <= spriteMemories_16_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1 <= spriteVisibleReg_16; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1 <= inSpriteHorizontal_16 & inSpriteVertical_16; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_16_REG <= spriteMemories_16_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_17_REG <= spriteMemories_17_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1 <= spriteVisibleReg_17; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1 <= inSpriteHorizontal_17 & inSpriteVertical_17; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_17_REG <= spriteMemories_17_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_18_REG <= spriteMemories_18_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1 <= spriteVisibleReg_18; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1 <= inSpriteHorizontal_18 & inSpriteVertical_18; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_18_REG <= spriteMemories_18_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_19_REG <= spriteMemories_19_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1 <= spriteVisibleReg_19; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1 <= inSpriteHorizontal_19 & inSpriteVertical_19; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_19_REG <= spriteMemories_19_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_20_REG <= spriteMemories_20_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1 <= spriteVisibleReg_20; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1 <= inSpriteHorizontal_20 & inSpriteVertical_20; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_20_REG <= spriteMemories_20_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_21_REG <= spriteMemories_21_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1 <= spriteVisibleReg_21; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1 <= inSpriteHorizontal_21 & inSpriteVertical_21; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_21_REG <= spriteMemories_21_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_22_REG <= spriteMemories_22_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1 <= spriteVisibleReg_22; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1 <= inSpriteHorizontal_22 & inSpriteVertical_22; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_22_REG <= spriteMemories_22_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_23_REG <= spriteMemories_23_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1 <= spriteVisibleReg_23; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1 <= inSpriteHorizontal_23 & inSpriteVertical_23; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_23_REG <= spriteMemories_23_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_24_REG <= spriteMemories_24_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1 <= spriteVisibleReg_24; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1 <= inSpriteHorizontal_24 & inSpriteVertical_24; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_24_REG <= spriteMemories_24_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_25_REG <= spriteMemories_25_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1 <= spriteVisibleReg_25; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1 <= inSpriteHorizontal_25 & inSpriteVertical_25; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_25_REG <= spriteMemories_25_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_26_REG <= spriteMemories_26_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1 <= spriteVisibleReg_26; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1 <= inSpriteHorizontal_26 & inSpriteVertical_26; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_26_REG <= spriteMemories_26_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_27_REG <= spriteMemories_27_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1 <= spriteVisibleReg_27; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1 <= inSpriteHorizontal_27 & inSpriteVertical_27; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_27_REG <= spriteMemories_27_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_28_REG <= spriteMemories_28_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1 <= spriteVisibleReg_28; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1 <= inSpriteHorizontal_28 & inSpriteVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_28_REG <= spriteMemories_28_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_29_REG <= spriteMemories_29_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1 <= spriteVisibleReg_29; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1 <= inSpriteHorizontal_28 & inSpriteVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_29_REG <= spriteMemories_29_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_30_REG <= spriteMemories_30_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1 <= spriteVisibleReg_30; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1 <= inSpriteHorizontal_28 & inSpriteVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_30_REG <= spriteMemories_30_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    multiHotPriortyReductionTree_io_dataInput_31_REG <= spriteMemories_31_io_dataRead[5:0]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 336:90]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 <=
      multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1 <= spriteVisibleReg_31; // @[\\src\\main\\scala\\GameUtilities.scala 23:30]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 <=
      multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1 <= inSpriteHorizontal_28 & inSpriteVertical_28; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 321:42]
    multiHotPriortyReductionTree_io_selectInput_31_REG <= spriteMemories_31_io_dataRead[6]; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 337:162]
    pixelColorSprite <= multiHotPriortyReductionTree_io_dataOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 339:33]
    pixelColorSpriteValid <= multiHotPriortyReductionTree_io_selectOutput; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 340:38]
    pixelColourVGA_pipeReg_0 <= pixelColourVGA_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    pixelColourVGA_pipeReg_1 <= pixelColourVGA_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 25:20]
    pixelColourVGA_pipeReg_2 <= CounterXReg < 10'h280 & CounterYReg < 10'h1e0; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 97:60]
    io_vgaRed_REG <= {pixelColourVGA[5:4],pixelColourVGA[5:4]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 346:26]
    io_vgaGreen_REG <= {pixelColourVGA[3:2],pixelColourVGA[3:2]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 347:28]
    io_vgaBlue_REG <= {pixelColourVGA[1:0],pixelColourVGA[1:0]}; // @[\\src\\main\\scala\\GraphicEngineVGA.scala 348:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ScaleCounterReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  CounterXReg = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  CounterYReg = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  backMemoryRestoreCounter = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  io_Hsync_pipeReg_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_Hsync_pipeReg_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_Hsync_pipeReg_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_Hsync_pipeReg_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_Vsync_pipeReg_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  io_Vsync_pipeReg_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_Vsync_pipeReg_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  io_Vsync_pipeReg_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  frameClockCount = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXPositionReg_0 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXPositionReg_1 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXPositionReg_2 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXPositionReg_3 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXPositionReg_4 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXPositionReg_5 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXPositionReg_6 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteXPositionReg_7 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  spriteXPositionReg_8 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  spriteXPositionReg_9 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  spriteXPositionReg_10 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  spriteXPositionReg_11 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  spriteXPositionReg_12 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  spriteXPositionReg_13 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  spriteXPositionReg_14 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  spriteXPositionReg_15 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  spriteXPositionReg_16 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  spriteXPositionReg_17 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  spriteXPositionReg_18 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  spriteXPositionReg_19 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  spriteXPositionReg_20 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  spriteXPositionReg_21 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  spriteXPositionReg_22 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  spriteXPositionReg_23 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  spriteXPositionReg_24 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  spriteXPositionReg_25 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  spriteXPositionReg_26 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  spriteXPositionReg_27 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  spriteYPositionReg_0 = _RAND_41[9:0];
  _RAND_42 = {1{`RANDOM}};
  spriteYPositionReg_1 = _RAND_42[9:0];
  _RAND_43 = {1{`RANDOM}};
  spriteYPositionReg_2 = _RAND_43[9:0];
  _RAND_44 = {1{`RANDOM}};
  spriteYPositionReg_3 = _RAND_44[9:0];
  _RAND_45 = {1{`RANDOM}};
  spriteYPositionReg_4 = _RAND_45[9:0];
  _RAND_46 = {1{`RANDOM}};
  spriteYPositionReg_5 = _RAND_46[9:0];
  _RAND_47 = {1{`RANDOM}};
  spriteYPositionReg_6 = _RAND_47[9:0];
  _RAND_48 = {1{`RANDOM}};
  spriteYPositionReg_7 = _RAND_48[9:0];
  _RAND_49 = {1{`RANDOM}};
  spriteYPositionReg_8 = _RAND_49[9:0];
  _RAND_50 = {1{`RANDOM}};
  spriteYPositionReg_9 = _RAND_50[9:0];
  _RAND_51 = {1{`RANDOM}};
  spriteYPositionReg_10 = _RAND_51[9:0];
  _RAND_52 = {1{`RANDOM}};
  spriteYPositionReg_11 = _RAND_52[9:0];
  _RAND_53 = {1{`RANDOM}};
  spriteYPositionReg_12 = _RAND_53[9:0];
  _RAND_54 = {1{`RANDOM}};
  spriteYPositionReg_13 = _RAND_54[9:0];
  _RAND_55 = {1{`RANDOM}};
  spriteYPositionReg_14 = _RAND_55[9:0];
  _RAND_56 = {1{`RANDOM}};
  spriteYPositionReg_15 = _RAND_56[9:0];
  _RAND_57 = {1{`RANDOM}};
  spriteYPositionReg_16 = _RAND_57[9:0];
  _RAND_58 = {1{`RANDOM}};
  spriteYPositionReg_17 = _RAND_58[9:0];
  _RAND_59 = {1{`RANDOM}};
  spriteYPositionReg_18 = _RAND_59[9:0];
  _RAND_60 = {1{`RANDOM}};
  spriteYPositionReg_19 = _RAND_60[9:0];
  _RAND_61 = {1{`RANDOM}};
  spriteYPositionReg_20 = _RAND_61[9:0];
  _RAND_62 = {1{`RANDOM}};
  spriteYPositionReg_21 = _RAND_62[9:0];
  _RAND_63 = {1{`RANDOM}};
  spriteYPositionReg_22 = _RAND_63[9:0];
  _RAND_64 = {1{`RANDOM}};
  spriteYPositionReg_23 = _RAND_64[9:0];
  _RAND_65 = {1{`RANDOM}};
  spriteYPositionReg_24 = _RAND_65[9:0];
  _RAND_66 = {1{`RANDOM}};
  spriteYPositionReg_25 = _RAND_66[9:0];
  _RAND_67 = {1{`RANDOM}};
  spriteYPositionReg_26 = _RAND_67[9:0];
  _RAND_68 = {1{`RANDOM}};
  spriteYPositionReg_27 = _RAND_68[9:0];
  _RAND_69 = {1{`RANDOM}};
  spriteVisibleReg_0 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  spriteVisibleReg_1 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  spriteVisibleReg_2 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  spriteVisibleReg_3 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  spriteVisibleReg_4 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  spriteVisibleReg_5 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  spriteVisibleReg_6 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  spriteVisibleReg_7 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  spriteVisibleReg_8 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  spriteVisibleReg_9 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  spriteVisibleReg_10 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  spriteVisibleReg_11 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  spriteVisibleReg_12 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  spriteVisibleReg_13 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  spriteVisibleReg_14 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  spriteVisibleReg_15 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  spriteVisibleReg_16 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  spriteVisibleReg_17 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  spriteVisibleReg_18 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  spriteVisibleReg_19 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  spriteVisibleReg_20 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  spriteVisibleReg_21 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  spriteVisibleReg_22 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  spriteVisibleReg_23 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  spriteVisibleReg_24 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  spriteVisibleReg_25 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  spriteVisibleReg_26 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  spriteVisibleReg_27 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  spriteVisibleReg_28 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  spriteVisibleReg_29 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  spriteVisibleReg_30 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  spriteVisibleReg_31 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  viewBoxXReg = _RAND_101[9:0];
  _RAND_102 = {1{`RANDOM}};
  viewBoxYReg = _RAND_102[8:0];
  _RAND_103 = {1{`RANDOM}};
  missingFrameErrorReg = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  backBufferWriteErrorReg = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  viewBoxOutOfRangeErrorReg = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  newFrameStikyReg = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  REG = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  backTileMemoryDataRead_0_REG = _RAND_108[6:0];
  _RAND_109 = {1{`RANDOM}};
  backTileMemoryDataRead_1_REG = _RAND_109[6:0];
  _RAND_110 = {1{`RANDOM}};
  backTileMemoryDataRead_2_REG = _RAND_110[6:0];
  _RAND_111 = {1{`RANDOM}};
  backTileMemoryDataRead_3_REG = _RAND_111[6:0];
  _RAND_112 = {1{`RANDOM}};
  backTileMemoryDataRead_4_REG = _RAND_112[6:0];
  _RAND_113 = {1{`RANDOM}};
  backTileMemoryDataRead_5_REG = _RAND_113[6:0];
  _RAND_114 = {1{`RANDOM}};
  backTileMemoryDataRead_6_REG = _RAND_114[6:0];
  _RAND_115 = {1{`RANDOM}};
  backTileMemoryDataRead_7_REG = _RAND_115[6:0];
  _RAND_116 = {1{`RANDOM}};
  backTileMemoryDataRead_8_REG = _RAND_116[6:0];
  _RAND_117 = {1{`RANDOM}};
  backTileMemoryDataRead_9_REG = _RAND_117[6:0];
  _RAND_118 = {1{`RANDOM}};
  backTileMemoryDataRead_10_REG = _RAND_118[6:0];
  _RAND_119 = {1{`RANDOM}};
  backTileMemoryDataRead_11_REG = _RAND_119[6:0];
  _RAND_120 = {1{`RANDOM}};
  backTileMemoryDataRead_12_REG = _RAND_120[6:0];
  _RAND_121 = {1{`RANDOM}};
  backTileMemoryDataRead_13_REG = _RAND_121[6:0];
  _RAND_122 = {1{`RANDOM}};
  backTileMemoryDataRead_14_REG = _RAND_122[6:0];
  _RAND_123 = {1{`RANDOM}};
  backTileMemoryDataRead_15_REG = _RAND_123[6:0];
  _RAND_124 = {1{`RANDOM}};
  backTileMemoryDataRead_16_REG = _RAND_124[6:0];
  _RAND_125 = {1{`RANDOM}};
  backTileMemoryDataRead_17_REG = _RAND_125[6:0];
  _RAND_126 = {1{`RANDOM}};
  backTileMemoryDataRead_18_REG = _RAND_126[6:0];
  _RAND_127 = {1{`RANDOM}};
  backTileMemoryDataRead_19_REG = _RAND_127[6:0];
  _RAND_128 = {1{`RANDOM}};
  backTileMemoryDataRead_20_REG = _RAND_128[6:0];
  _RAND_129 = {1{`RANDOM}};
  backTileMemoryDataRead_21_REG = _RAND_129[6:0];
  _RAND_130 = {1{`RANDOM}};
  backTileMemoryDataRead_22_REG = _RAND_130[6:0];
  _RAND_131 = {1{`RANDOM}};
  backTileMemoryDataRead_23_REG = _RAND_131[6:0];
  _RAND_132 = {1{`RANDOM}};
  backTileMemoryDataRead_24_REG = _RAND_132[6:0];
  _RAND_133 = {1{`RANDOM}};
  backTileMemoryDataRead_25_REG = _RAND_133[6:0];
  _RAND_134 = {1{`RANDOM}};
  backTileMemoryDataRead_26_REG = _RAND_134[6:0];
  _RAND_135 = {1{`RANDOM}};
  backTileMemoryDataRead_27_REG = _RAND_135[6:0];
  _RAND_136 = {1{`RANDOM}};
  backTileMemoryDataRead_28_REG = _RAND_136[6:0];
  _RAND_137 = {1{`RANDOM}};
  backTileMemoryDataRead_29_REG = _RAND_137[6:0];
  _RAND_138 = {1{`RANDOM}};
  backTileMemoryDataRead_30_REG = _RAND_138[6:0];
  _RAND_139 = {1{`RANDOM}};
  backTileMemoryDataRead_31_REG = _RAND_139[6:0];
  _RAND_140 = {1{`RANDOM}};
  backMemoryCopyCounter = _RAND_140[11:0];
  _RAND_141 = {1{`RANDOM}};
  copyEnabledReg = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  backBufferShadowMemory_io_address_REG = _RAND_142[10:0];
  _RAND_143 = {1{`RANDOM}};
  backBufferShadowMemory_io_address_REG_1 = _RAND_143[10:0];
  _RAND_144 = {1{`RANDOM}};
  backBufferShadowMemory_io_writeEnable_REG = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  backBufferShadowMemory_io_writeEnable_REG_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  backBufferShadowMemory_io_dataWrite_REG = _RAND_146[4:0];
  _RAND_147 = {1{`RANDOM}};
  backBufferMemory_io_address_REG = _RAND_147[10:0];
  _RAND_148 = {1{`RANDOM}};
  fullBackgroundColor_REG = _RAND_148[4:0];
  _RAND_149 = {1{`RANDOM}};
  pixelColorBack = _RAND_149[5:0];
  _RAND_150 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_0_REG = _RAND_150[5:0];
  _RAND_151 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg__1 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_0 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_pipeReg_1_1 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_0_REG = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_1_REG = _RAND_156[5:0];
  _RAND_157 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg__1 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_0 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_pipeReg_1_1 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_1_REG = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_2_REG = _RAND_162[5:0];
  _RAND_163 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg__1 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_0 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_pipeReg_1_1 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_2_REG = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_3_REG = _RAND_168[5:0];
  _RAND_169 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg__1 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_0 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_pipeReg_1_1 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_3_REG = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_4_REG = _RAND_174[5:0];
  _RAND_175 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg__1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_0 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_pipeReg_1_1 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_4_REG = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_5_REG = _RAND_180[5:0];
  _RAND_181 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg__1 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_pipeReg_1_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_5_REG = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_6_REG = _RAND_186[5:0];
  _RAND_187 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg__1 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_0 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_pipeReg_1_1 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_6_REG = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_7_REG = _RAND_192[5:0];
  _RAND_193 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__0 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg__1 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_0 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_pipeReg_1_1 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_7_REG = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_8_REG = _RAND_198[5:0];
  _RAND_199 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg__1 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_0 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_pipeReg_1_1 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_8_REG = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_9_REG = _RAND_204[5:0];
  _RAND_205 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg__1 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_0 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_pipeReg_1_1 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_9_REG = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_10_REG = _RAND_210[5:0];
  _RAND_211 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg__1 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_0 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_pipeReg_1_1 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_10_REG = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_11_REG = _RAND_216[5:0];
  _RAND_217 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__0 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg__1 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_0 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_pipeReg_1_1 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_11_REG = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_12_REG = _RAND_222[5:0];
  _RAND_223 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg__1 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_0 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_pipeReg_1_1 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_12_REG = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_13_REG = _RAND_228[5:0];
  _RAND_229 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__0 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg__1 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_0 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_pipeReg_1_1 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_13_REG = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_14_REG = _RAND_234[5:0];
  _RAND_235 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg__1 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_0 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_pipeReg_1_1 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_14_REG = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_15_REG = _RAND_240[5:0];
  _RAND_241 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg__1 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_0 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_pipeReg_1_1 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_15_REG = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_16_REG = _RAND_246[5:0];
  _RAND_247 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg__1 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_0 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_pipeReg_1_1 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_16_REG = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_17_REG = _RAND_252[5:0];
  _RAND_253 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__0 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg__1 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_0 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_pipeReg_1_1 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_17_REG = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_18_REG = _RAND_258[5:0];
  _RAND_259 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg__1 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_0 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_pipeReg_1_1 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_18_REG = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_19_REG = _RAND_264[5:0];
  _RAND_265 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__0 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg__1 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_0 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_pipeReg_1_1 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_19_REG = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_20_REG = _RAND_270[5:0];
  _RAND_271 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__0 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg__1 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_0 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_pipeReg_1_1 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_20_REG = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_21_REG = _RAND_276[5:0];
  _RAND_277 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__0 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg__1 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_0 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_pipeReg_1_1 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_21_REG = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_22_REG = _RAND_282[5:0];
  _RAND_283 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg__1 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_0 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_pipeReg_1_1 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_22_REG = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_23_REG = _RAND_288[5:0];
  _RAND_289 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__0 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg__1 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_0 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_pipeReg_1_1 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_23_REG = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_24_REG = _RAND_294[5:0];
  _RAND_295 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__0 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg__1 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_0 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_pipeReg_1_1 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_24_REG = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_25_REG = _RAND_300[5:0];
  _RAND_301 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__0 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg__1 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_0 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_pipeReg_1_1 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_25_REG = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_26_REG = _RAND_306[5:0];
  _RAND_307 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg__1 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_0 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_pipeReg_1_1 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_26_REG = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_27_REG = _RAND_312[5:0];
  _RAND_313 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__0 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg__1 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_0 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_pipeReg_1_1 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_27_REG = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_28_REG = _RAND_318[5:0];
  _RAND_319 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__0 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg__1 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_0 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_pipeReg_1_1 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_28_REG = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_29_REG = _RAND_324[5:0];
  _RAND_325 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__0 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg__1 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_0 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_pipeReg_1_1 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_29_REG = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_30_REG = _RAND_330[5:0];
  _RAND_331 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__0 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg__1 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_0 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_pipeReg_1_1 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_30_REG = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_dataInput_31_REG = _RAND_336[5:0];
  _RAND_337 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg__1 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_0 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_pipeReg_1_1 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  multiHotPriortyReductionTree_io_selectInput_31_REG = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  pixelColorSprite = _RAND_342[5:0];
  _RAND_343 = {1{`RANDOM}};
  pixelColorSpriteValid = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_0 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  pixelColourVGA_pipeReg_2 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  io_vgaRed_REG = _RAND_347[3:0];
  _RAND_348 = {1{`RANDOM}};
  io_vgaGreen_REG = _RAND_348[3:0];
  _RAND_349 = {1{`RANDOM}};
  io_vgaBlue_REG = _RAND_349[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Memory_67(
  input         clock,
  input  [7:0]  io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [27:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [7:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(8), .DATA_WIDTH(28), .LOAD_FILE("memory_init/tune_init_0.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 28'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module Memory_68(
  input         clock,
  input  [7:0]  io_address, // @[\\src\\main\\scala\\Memory.scala 48:14]
  output [27:0] io_dataRead // @[\\src\\main\\scala\\Memory.scala 48:14]
);
  wire  ramsSpWf_clk; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_we; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire  ramsSpWf_en; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [7:0] ramsSpWf_addr; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_di; // @[\\src\\main\\scala\\Memory.scala 65:26]
  wire [27:0] ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(8), .DATA_WIDTH(28), .LOAD_FILE("memory_init/tune_init_1.mem")) ramsSpWf ( // @[\\src\\main\\scala\\Memory.scala 65:26]
    .clk(ramsSpWf_clk),
    .we(ramsSpWf_we),
    .en(ramsSpWf_en),
    .addr(ramsSpWf_addr),
    .di(ramsSpWf_di),
    .dout(ramsSpWf_dout)
  );
  assign io_dataRead = ramsSpWf_dout; // @[\\src\\main\\scala\\Memory.scala 71:17]
  assign ramsSpWf_clk = clock; // @[\\src\\main\\scala\\Memory.scala 66:21]
  assign ramsSpWf_we = 1'h0; // @[\\src\\main\\scala\\Memory.scala 67:20]
  assign ramsSpWf_en = 1'h1; // @[\\src\\main\\scala\\Memory.scala 68:20]
  assign ramsSpWf_addr = io_address; // @[\\src\\main\\scala\\Memory.scala 69:22]
  assign ramsSpWf_di = 28'h0; // @[\\src\\main\\scala\\Memory.scala 70:20]
endmodule
module SoundEngine(
  input   clock,
  input   reset,
  output  io_soundOut, // @[\\src\\main\\scala\\SoundEngine.scala 13:14]
  input   io_startTune_0 // @[\\src\\main\\scala\\SoundEngine.scala 13:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  tuneMemories_0_clock; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [7:0] tuneMemories_0_io_address; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [27:0] tuneMemories_0_io_dataRead; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire  tuneMemories_1_clock; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [7:0] tuneMemories_1_io_address; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  wire [27:0] tuneMemories_1_io_dataRead; // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
  reg [16:0] counter1msReg; // @[\\src\\main\\scala\\SoundEngine.scala 34:30]
  wire  enable1ms = counter1msReg == 17'h0; // @[\\src\\main\\scala\\SoundEngine.scala 35:33]
  wire [16:0] _counter1msReg_T_2 = counter1msReg - 17'h1; // @[\\src\\main\\scala\\SoundEngine.scala 36:90]
  reg [4:0] counter32ccReg; // @[\\src\\main\\scala\\SoundEngine.scala 38:31]
  wire  enable32cc = counter32ccReg == 5'h0; // @[\\src\\main\\scala\\SoundEngine.scala 39:35]
  wire [4:0] _counter32ccReg_T_2 = counter32ccReg - 5'h1; // @[\\src\\main\\scala\\SoundEngine.scala 40:95]
  reg [15:0] noteCountReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 44:29]
  reg [11:0] durationCountReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
  reg [11:0] durationCountReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
  reg [15:0] currNoteReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 57:28]
  reg [11:0] currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
  reg [11:0] currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
  reg [7:0] nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
  reg [7:0] nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
  reg [1:0] stateReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
  reg [1:0] stateReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
  reg  newNoteLoadReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
  reg  newNoteLoadReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
  reg  audioReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 64:25]
  reg  isPlayingReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 65:29]
  wire  noteCountRegEnable_0 = isPlayingReg_0 & enable32cc; // @[\\src\\main\\scala\\SoundEngine.scala 74:46]
  wire  durationCountRegEnable_0 = isPlayingReg_0 & enable1ms; // @[\\src\\main\\scala\\SoundEngine.scala 75:50]
  wire [15:0] _noteCountReg_0_T_1 = noteCountReg_0 - 16'h1; // @[\\src\\main\\scala\\SoundEngine.scala 80:42]
  wire  noteCountRegDone_0 = noteCountReg_0 == 16'h0; // @[\\src\\main\\scala\\SoundEngine.scala 82:46]
  wire  noteCountRegLoad_0 = noteCountRegDone_0 | newNoteLoadReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 91:48]
  wire [11:0] _durationCountReg_0_T_1 = durationCountReg_0 - 12'h1; // @[\\src\\main\\scala\\SoundEngine.scala 87:50]
  wire  durationCountRegDone_0 = durationCountReg_0 == 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 89:54]
  wire  _T_8 = tuneMemories_0_io_dataRead[27:16] != 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 111:60]
  wire [1:0] _GEN_4 = tuneMemories_0_io_dataRead[27:16] != 12'h0 ? 2'h3 : stateReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 112:23 62:25]
  wire [15:0] _GEN_5 = tuneMemories_0_io_dataRead[27:16] != 12'h0 ? tuneMemories_0_io_dataRead[15:0] : currNoteReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 113:26 57:28]
  wire [11:0] _GEN_6 = tuneMemories_0_io_dataRead[27:16] != 12'h0 ? tuneMemories_0_io_dataRead[27:16] :
    currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 114:30 58:32]
  wire  _T_13 = durationCountRegDone_0 & ~newNoteLoadReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:44]
  wire [7:0] _nextIndexReg_0_T_1 = nextIndexReg_0 + 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 126:46]
  wire  _GEN_8 = nextIndexReg_0 == 8'h0 ? 1'h0 : isPlayingReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 127:40 128:29 65:29]
  wire [15:0] _GEN_9 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? tuneMemories_0_io_dataRead[15:0] : currNoteReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 123:26 57:28]
  wire [11:0] _GEN_10 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? tuneMemories_0_io_dataRead[27:16] :
    currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 124:30 58:32]
  wire [7:0] _GEN_12 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? _nextIndexReg_0_T_1 : nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 126:27 59:29]
  wire  _GEN_13 = durationCountRegDone_0 & ~newNoteLoadReg_0 ? _GEN_8 : isPlayingReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 65:29]
  wire [7:0] _GEN_14 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? 8'h0 : _GEN_12; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 120:27]
  wire [15:0] _GEN_15 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? currNoteReg_0 : _GEN_9; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 57:28]
  wire [11:0] _GEN_16 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? currDurationReg_0 : _GEN_10; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 58:32]
  wire  _GEN_17 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? 1'h0 : _T_13; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 97:23]
  wire  _GEN_18 = tuneMemories_0_io_dataRead[27:16] == 12'h0 ? isPlayingReg_0 : _GEN_13; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 65:29]
  wire  _GEN_20 = io_startTune_0 | _GEN_18; // @[\\src\\main\\scala\\SoundEngine.scala 134:32 135:27]
  wire [7:0] _GEN_22 = 2'h3 == stateReg_0 ? _GEN_14 : nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 59:29]
  wire [15:0] _GEN_23 = 2'h3 == stateReg_0 ? _GEN_15 : currNoteReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 57:28]
  wire [11:0] _GEN_24 = 2'h3 == stateReg_0 ? _GEN_16 : currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 58:32]
  wire  _GEN_25 = 2'h3 == stateReg_0 & _GEN_17; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 97:23]
  wire  _GEN_26 = 2'h3 == stateReg_0 ? _GEN_20 : isPlayingReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 65:29]
  wire  _GEN_46 = noteCountRegDone_0 ? ~audioReg_0 : audioReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 145:33 146:21 64:25]
  wire  _GEN_47 = isPlayingReg_0 & currNoteReg_0 != 16'h0 & _GEN_46; // @[\\src\\main\\scala\\SoundEngine.scala 144:53 149:19]
  wire  durationCountRegDone_1 = durationCountReg_1 == 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 89:54]
  wire  _T_25 = tuneMemories_1_io_dataRead[27:16] != 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 111:60]
  wire [1:0] _GEN_52 = tuneMemories_1_io_dataRead[27:16] != 12'h0 ? 2'h3 : stateReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 112:23 62:25]
  wire [11:0] _GEN_54 = tuneMemories_1_io_dataRead[27:16] != 12'h0 ? tuneMemories_1_io_dataRead[27:16] :
    currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 111:69 114:30 58:32]
  wire  _T_30 = durationCountRegDone_1 & ~newNoteLoadReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:44]
  wire [7:0] _nextIndexReg_1_T_1 = nextIndexReg_1 + 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 126:46]
  wire [11:0] _GEN_58 = durationCountRegDone_1 & ~newNoteLoadReg_1 ? tuneMemories_1_io_dataRead[27:16] :
    currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 124:30 58:32]
  wire [7:0] _GEN_60 = durationCountRegDone_1 & ~newNoteLoadReg_1 ? _nextIndexReg_1_T_1 : nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 122:67 126:27 59:29]
  wire [7:0] _GEN_62 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? 8'h0 : _GEN_60; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 120:27]
  wire [11:0] _GEN_64 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? currDurationReg_1 : _GEN_58; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 58:32]
  wire  _GEN_65 = tuneMemories_1_io_dataRead[27:16] == 12'h0 ? 1'h0 : _T_30; // @[\\src\\main\\scala\\SoundEngine.scala 119:69 97:23]
  wire [7:0] _GEN_70 = 2'h3 == stateReg_1 ? _GEN_62 : nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 59:29]
  wire [11:0] _GEN_72 = 2'h3 == stateReg_1 ? _GEN_64 : currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 58:32]
  wire  _GEN_73 = 2'h3 == stateReg_1 & _GEN_65; // @[\\src\\main\\scala\\SoundEngine.scala 100:25 97:23]
  Memory_67 tuneMemories_0 ( // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
    .clock(tuneMemories_0_clock),
    .io_address(tuneMemories_0_io_address),
    .io_dataRead(tuneMemories_0_io_dataRead)
  );
  Memory_68 tuneMemories_1 ( // @[\\src\\main\\scala\\SoundEngine.scala 26:28]
    .clock(tuneMemories_1_clock),
    .io_address(tuneMemories_1_io_address),
    .io_dataRead(tuneMemories_1_io_dataRead)
  );
  assign io_soundOut = audioReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 155:{15,15}]
  assign tuneMemories_0_clock = clock;
  assign tuneMemories_0_io_address = nextIndexReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 72:32]
  assign tuneMemories_1_clock = clock;
  assign tuneMemories_1_io_address = nextIndexReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 72:32]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 34:30]
      counter1msReg <= 17'h1869f; // @[\\src\\main\\scala\\SoundEngine.scala 34:30]
    end else if (enable1ms) begin // @[\\src\\main\\scala\\SoundEngine.scala 36:23]
      counter1msReg <= 17'h1869f;
    end else begin
      counter1msReg <= _counter1msReg_T_2;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 38:31]
      counter32ccReg <= 5'h1f; // @[\\src\\main\\scala\\SoundEngine.scala 38:31]
    end else if (enable32cc) begin // @[\\src\\main\\scala\\SoundEngine.scala 40:24]
      counter32ccReg <= 5'h1f;
    end else begin
      counter32ccReg <= _counter32ccReg_T_2;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 44:29]
      noteCountReg_0 <= 16'h0; // @[\\src\\main\\scala\\SoundEngine.scala 44:29]
    end else if (noteCountRegLoad_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 77:31]
      noteCountReg_0 <= currNoteReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 78:23]
    end else if (noteCountRegEnable_0 & noteCountReg_0 != 16'h0) begin // @[\\src\\main\\scala\\SoundEngine.scala 79:66]
      noteCountReg_0 <= _noteCountReg_0_T_1; // @[\\src\\main\\scala\\SoundEngine.scala 80:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
      durationCountReg_0 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
    end else if (newNoteLoadReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 84:35]
      durationCountReg_0 <= currDurationReg_0; // @[\\src\\main\\scala\\SoundEngine.scala 85:27]
    end else if (durationCountRegEnable_0 & durationCountReg_0 != 12'h0) begin // @[\\src\\main\\scala\\SoundEngine.scala 86:74]
      durationCountReg_0 <= _durationCountReg_0_T_1; // @[\\src\\main\\scala\\SoundEngine.scala 87:27]
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
      durationCountReg_1 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 45:33]
    end else if (newNoteLoadReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 84:35]
      durationCountReg_1 <= currDurationReg_1; // @[\\src\\main\\scala\\SoundEngine.scala 85:27]
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 57:28]
      currNoteReg_0 <= 16'h0; // @[\\src\\main\\scala\\SoundEngine.scala 57:28]
    end else if (!(2'h0 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h1 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
          currNoteReg_0 <= _GEN_5;
        end else begin
          currNoteReg_0 <= _GEN_23;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
      currDurationReg_0 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
    end else if (!(2'h0 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h1 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
          currDurationReg_0 <= _GEN_6;
        end else begin
          currDurationReg_0 <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
      currDurationReg_1 <= 12'h0; // @[\\src\\main\\scala\\SoundEngine.scala 58:32]
    end else if (!(2'h0 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h1 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
          currDurationReg_1 <= _GEN_54;
        end else begin
          currDurationReg_1 <= _GEN_72;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
      nextIndexReg_0 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 102:25]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 107:25]
    end else if (!(2'h2 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_0 <= _GEN_22;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
      nextIndexReg_1 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 59:29]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= 8'h0; // @[\\src\\main\\scala\\SoundEngine.scala 102:25]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= 8'h1; // @[\\src\\main\\scala\\SoundEngine.scala 107:25]
    end else if (!(2'h2 == stateReg_1)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      nextIndexReg_1 <= _GEN_70;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
      stateReg_0 <= 2'h0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= 2'h1; // @[\\src\\main\\scala\\SoundEngine.scala 103:21]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= 2'h2; // @[\\src\\main\\scala\\SoundEngine.scala 108:21]
    end else if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_0 <= _GEN_4;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
      stateReg_1 <= 2'h0; // @[\\src\\main\\scala\\SoundEngine.scala 62:25]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= 2'h1; // @[\\src\\main\\scala\\SoundEngine.scala 103:21]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= 2'h2; // @[\\src\\main\\scala\\SoundEngine.scala 108:21]
    end else if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      stateReg_1 <= _GEN_52;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h1 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h2 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_0 <= _T_8;
    end else begin
      newNoteLoadReg_0 <= _GEN_25;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 63:31]
    end else if (2'h0 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h1 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 97:23]
    end else if (2'h2 == stateReg_1) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      newNoteLoadReg_1 <= _T_25;
    end else begin
      newNoteLoadReg_1 <= _GEN_73;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 64:25]
      audioReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 64:25]
    end else begin
      audioReg_0 <= _GEN_47;
    end
    if (reset) begin // @[\\src\\main\\scala\\SoundEngine.scala 65:29]
      isPlayingReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 65:29]
    end else if (2'h0 == stateReg_0) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      isPlayingReg_0 <= 1'h0; // @[\\src\\main\\scala\\SoundEngine.scala 104:25]
    end else if (!(2'h1 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
      if (!(2'h2 == stateReg_0)) begin // @[\\src\\main\\scala\\SoundEngine.scala 100:25]
        isPlayingReg_0 <= _GEN_26;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter1msReg = _RAND_0[16:0];
  _RAND_1 = {1{`RANDOM}};
  counter32ccReg = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  noteCountReg_0 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  durationCountReg_0 = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  durationCountReg_1 = _RAND_4[11:0];
  _RAND_5 = {1{`RANDOM}};
  currNoteReg_0 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  currDurationReg_0 = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  currDurationReg_1 = _RAND_7[11:0];
  _RAND_8 = {1{`RANDOM}};
  nextIndexReg_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  nextIndexReg_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  stateReg_0 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  stateReg_1 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  newNoteLoadReg_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  newNoteLoadReg_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  audioReg_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  isPlayingReg_0 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PosToGridIndex(
  input  [10:0] io_xPos, // @[\\src\\main\\scala\\PosToGridIndex.scala 12:14]
  input  [9:0]  io_yPos, // @[\\src\\main\\scala\\PosToGridIndex.scala 12:14]
  output [8:0]  io_index // @[\\src\\main\\scala\\PosToGridIndex.scala 12:14]
);
  wire [9:0] _io_index_T_3 = $signed(io_yPos) - 10'sh4; // @[\\src\\main\\scala\\PosToGridIndex.scala 18:31]
  wire [14:0] _io_index_T_4 = _io_index_T_3 * 5'h19; // @[\\src\\main\\scala\\PosToGridIndex.scala 18:38]
  wire [10:0] _io_index_T_8 = $signed(io_xPos) + 11'sh4; // @[\\src\\main\\scala\\PosToGridIndex.scala 18:63]
  wire [14:0] _GEN_0 = {{4'd0}, _io_index_T_8}; // @[\\src\\main\\scala\\PosToGridIndex.scala 18:45]
  wire [14:0] _io_index_T_10 = _io_index_T_4 + _GEN_0; // @[\\src\\main\\scala\\PosToGridIndex.scala 18:45]
  assign io_index = _io_index_T_10[8:0]; // @[\\src\\main\\scala\\PosToGridIndex.scala 18:12]
endmodule
module CollisionDetector(
  input  [2:0]  io_grid_0, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_1, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_2, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_3, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_4, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_5, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_6, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_7, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_8, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_9, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_10, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_11, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_12, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_13, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_14, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_15, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_16, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_17, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_18, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_19, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_20, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_21, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_22, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_23, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_24, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_25, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_26, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_27, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_28, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_29, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_30, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_31, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_32, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_33, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_34, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_35, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_36, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_37, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_38, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_39, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_40, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_41, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_42, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_43, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_44, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_45, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_46, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_47, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_48, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_49, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_50, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_51, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_52, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_53, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_54, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_55, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_56, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_57, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_58, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_59, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_60, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_61, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_62, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_63, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_64, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_65, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_66, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_67, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_68, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_69, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_70, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_71, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_72, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_73, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_74, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_75, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_76, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_77, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_78, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_79, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_80, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_81, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_82, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_83, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_84, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_85, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_86, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_87, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_88, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_89, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_90, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_91, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_92, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_93, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_94, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_95, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_96, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_97, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_98, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_99, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_100, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_101, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_102, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_103, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_104, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_105, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_106, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_107, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_108, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_109, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_110, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_111, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_112, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_113, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_114, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_115, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_116, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_117, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_118, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_119, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_120, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_121, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_122, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_123, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_124, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_125, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_126, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_127, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_128, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_129, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_130, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_131, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_132, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_133, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_134, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_135, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_136, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_137, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_138, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_139, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_140, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_141, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_142, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_143, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_144, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_145, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_146, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_147, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_148, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_149, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_150, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_151, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_152, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_153, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_154, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_155, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_156, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_157, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_158, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_159, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_160, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_161, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_162, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_163, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_164, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_165, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_166, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_167, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_168, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_169, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_170, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_171, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_172, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_173, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_174, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_175, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_176, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_177, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_178, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_179, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_180, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_181, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_182, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_183, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_184, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_185, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_186, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_187, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_188, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_189, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_190, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_191, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_192, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_193, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_194, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_195, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_196, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_197, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_198, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_199, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_200, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_201, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_202, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_203, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_204, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_205, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_206, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_207, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_208, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_209, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_210, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_211, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_212, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_213, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_214, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_215, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_216, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_217, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_218, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_219, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_220, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_221, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_222, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_223, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_224, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_225, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_226, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_227, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_228, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_229, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_230, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_231, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_232, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_233, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_234, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_235, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_236, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_237, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_238, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_239, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_240, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_241, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_242, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_243, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_244, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_245, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_246, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_247, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_248, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_249, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_250, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_251, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_252, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_253, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_254, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_255, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_256, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_257, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_258, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_259, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_260, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_261, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_262, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_263, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_264, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_265, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_266, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_267, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_268, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_269, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_270, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_271, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_272, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_273, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_274, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_275, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_276, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_277, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_278, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_279, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_280, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_281, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_282, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_283, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_284, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_285, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_286, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_287, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_288, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_289, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_290, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_291, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_292, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_293, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_294, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_295, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_296, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_297, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_298, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [2:0]  io_grid_299, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [10:0] io_xPos, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [9:0]  io_yPos, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [3:0]  io_xOffsets_0, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [3:0]  io_xOffsets_1, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [3:0]  io_xOffsets_2, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [3:0]  io_xOffsets_3, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [3:0]  io_yOffsets_0, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [3:0]  io_yOffsets_1, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [3:0]  io_yOffsets_2, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  input  [3:0]  io_yOffsets_3, // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
  output        io_isCollision // @[\\src\\main\\scala\\CollisionDetector.scala 12:14]
);
  wire [10:0] first_io_xPos; // @[\\src\\main\\scala\\CollisionDetector.scala 22:21]
  wire [9:0] first_io_yPos; // @[\\src\\main\\scala\\CollisionDetector.scala 22:21]
  wire [8:0] first_io_index; // @[\\src\\main\\scala\\CollisionDetector.scala 22:21]
  wire [10:0] second_io_xPos; // @[\\src\\main\\scala\\CollisionDetector.scala 23:22]
  wire [9:0] second_io_yPos; // @[\\src\\main\\scala\\CollisionDetector.scala 23:22]
  wire [8:0] second_io_index; // @[\\src\\main\\scala\\CollisionDetector.scala 23:22]
  wire [10:0] third_io_xPos; // @[\\src\\main\\scala\\CollisionDetector.scala 24:21]
  wire [9:0] third_io_yPos; // @[\\src\\main\\scala\\CollisionDetector.scala 24:21]
  wire [8:0] third_io_index; // @[\\src\\main\\scala\\CollisionDetector.scala 24:21]
  wire [10:0] fourth_io_xPos; // @[\\src\\main\\scala\\CollisionDetector.scala 25:23]
  wire [9:0] fourth_io_yPos; // @[\\src\\main\\scala\\CollisionDetector.scala 25:23]
  wire [8:0] fourth_io_index; // @[\\src\\main\\scala\\CollisionDetector.scala 25:23]
  wire [10:0] _GEN_1200 = {{7{io_xOffsets_0[3]}},io_xOffsets_0}; // @[\\src\\main\\scala\\CollisionDetector.scala 26:28]
  wire [9:0] _GEN_1201 = {{6{io_yOffsets_0[3]}},io_yOffsets_0}; // @[\\src\\main\\scala\\CollisionDetector.scala 27:28]
  wire [10:0] _GEN_1202 = {{7{io_xOffsets_1[3]}},io_xOffsets_1}; // @[\\src\\main\\scala\\CollisionDetector.scala 28:29]
  wire [9:0] _GEN_1203 = {{6{io_yOffsets_1[3]}},io_yOffsets_1}; // @[\\src\\main\\scala\\CollisionDetector.scala 29:29]
  wire [10:0] _GEN_1204 = {{7{io_xOffsets_2[3]}},io_xOffsets_2}; // @[\\src\\main\\scala\\CollisionDetector.scala 30:28]
  wire [9:0] _GEN_1205 = {{6{io_yOffsets_2[3]}},io_yOffsets_2}; // @[\\src\\main\\scala\\CollisionDetector.scala 31:28]
  wire [10:0] _GEN_1206 = {{7{io_xOffsets_3[3]}},io_xOffsets_3}; // @[\\src\\main\\scala\\CollisionDetector.scala 32:29]
  wire [9:0] _GEN_1207 = {{6{io_yOffsets_3[3]}},io_yOffsets_3}; // @[\\src\\main\\scala\\CollisionDetector.scala 33:29]
  wire [2:0] _GEN_1 = 9'h1 == first_io_index ? io_grid_1 : io_grid_0; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_2 = 9'h2 == first_io_index ? io_grid_2 : _GEN_1; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_3 = 9'h3 == first_io_index ? io_grid_3 : _GEN_2; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_4 = 9'h4 == first_io_index ? io_grid_4 : _GEN_3; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_5 = 9'h5 == first_io_index ? io_grid_5 : _GEN_4; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_6 = 9'h6 == first_io_index ? io_grid_6 : _GEN_5; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_7 = 9'h7 == first_io_index ? io_grid_7 : _GEN_6; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_8 = 9'h8 == first_io_index ? io_grid_8 : _GEN_7; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_9 = 9'h9 == first_io_index ? io_grid_9 : _GEN_8; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_10 = 9'ha == first_io_index ? io_grid_10 : _GEN_9; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_11 = 9'hb == first_io_index ? io_grid_11 : _GEN_10; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_12 = 9'hc == first_io_index ? io_grid_12 : _GEN_11; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_13 = 9'hd == first_io_index ? io_grid_13 : _GEN_12; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_14 = 9'he == first_io_index ? io_grid_14 : _GEN_13; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_15 = 9'hf == first_io_index ? io_grid_15 : _GEN_14; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_16 = 9'h10 == first_io_index ? io_grid_16 : _GEN_15; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_17 = 9'h11 == first_io_index ? io_grid_17 : _GEN_16; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_18 = 9'h12 == first_io_index ? io_grid_18 : _GEN_17; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_19 = 9'h13 == first_io_index ? io_grid_19 : _GEN_18; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_20 = 9'h14 == first_io_index ? io_grid_20 : _GEN_19; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_21 = 9'h15 == first_io_index ? io_grid_21 : _GEN_20; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_22 = 9'h16 == first_io_index ? io_grid_22 : _GEN_21; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_23 = 9'h17 == first_io_index ? io_grid_23 : _GEN_22; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_24 = 9'h18 == first_io_index ? io_grid_24 : _GEN_23; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_25 = 9'h19 == first_io_index ? io_grid_25 : _GEN_24; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_26 = 9'h1a == first_io_index ? io_grid_26 : _GEN_25; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_27 = 9'h1b == first_io_index ? io_grid_27 : _GEN_26; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_28 = 9'h1c == first_io_index ? io_grid_28 : _GEN_27; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_29 = 9'h1d == first_io_index ? io_grid_29 : _GEN_28; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_30 = 9'h1e == first_io_index ? io_grid_30 : _GEN_29; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_31 = 9'h1f == first_io_index ? io_grid_31 : _GEN_30; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_32 = 9'h20 == first_io_index ? io_grid_32 : _GEN_31; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_33 = 9'h21 == first_io_index ? io_grid_33 : _GEN_32; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_34 = 9'h22 == first_io_index ? io_grid_34 : _GEN_33; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_35 = 9'h23 == first_io_index ? io_grid_35 : _GEN_34; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_36 = 9'h24 == first_io_index ? io_grid_36 : _GEN_35; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_37 = 9'h25 == first_io_index ? io_grid_37 : _GEN_36; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_38 = 9'h26 == first_io_index ? io_grid_38 : _GEN_37; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_39 = 9'h27 == first_io_index ? io_grid_39 : _GEN_38; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_40 = 9'h28 == first_io_index ? io_grid_40 : _GEN_39; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_41 = 9'h29 == first_io_index ? io_grid_41 : _GEN_40; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_42 = 9'h2a == first_io_index ? io_grid_42 : _GEN_41; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_43 = 9'h2b == first_io_index ? io_grid_43 : _GEN_42; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_44 = 9'h2c == first_io_index ? io_grid_44 : _GEN_43; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_45 = 9'h2d == first_io_index ? io_grid_45 : _GEN_44; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_46 = 9'h2e == first_io_index ? io_grid_46 : _GEN_45; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_47 = 9'h2f == first_io_index ? io_grid_47 : _GEN_46; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_48 = 9'h30 == first_io_index ? io_grid_48 : _GEN_47; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_49 = 9'h31 == first_io_index ? io_grid_49 : _GEN_48; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_50 = 9'h32 == first_io_index ? io_grid_50 : _GEN_49; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_51 = 9'h33 == first_io_index ? io_grid_51 : _GEN_50; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_52 = 9'h34 == first_io_index ? io_grid_52 : _GEN_51; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_53 = 9'h35 == first_io_index ? io_grid_53 : _GEN_52; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_54 = 9'h36 == first_io_index ? io_grid_54 : _GEN_53; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_55 = 9'h37 == first_io_index ? io_grid_55 : _GEN_54; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_56 = 9'h38 == first_io_index ? io_grid_56 : _GEN_55; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_57 = 9'h39 == first_io_index ? io_grid_57 : _GEN_56; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_58 = 9'h3a == first_io_index ? io_grid_58 : _GEN_57; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_59 = 9'h3b == first_io_index ? io_grid_59 : _GEN_58; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_60 = 9'h3c == first_io_index ? io_grid_60 : _GEN_59; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_61 = 9'h3d == first_io_index ? io_grid_61 : _GEN_60; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_62 = 9'h3e == first_io_index ? io_grid_62 : _GEN_61; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_63 = 9'h3f == first_io_index ? io_grid_63 : _GEN_62; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_64 = 9'h40 == first_io_index ? io_grid_64 : _GEN_63; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_65 = 9'h41 == first_io_index ? io_grid_65 : _GEN_64; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_66 = 9'h42 == first_io_index ? io_grid_66 : _GEN_65; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_67 = 9'h43 == first_io_index ? io_grid_67 : _GEN_66; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_68 = 9'h44 == first_io_index ? io_grid_68 : _GEN_67; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_69 = 9'h45 == first_io_index ? io_grid_69 : _GEN_68; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_70 = 9'h46 == first_io_index ? io_grid_70 : _GEN_69; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_71 = 9'h47 == first_io_index ? io_grid_71 : _GEN_70; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_72 = 9'h48 == first_io_index ? io_grid_72 : _GEN_71; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_73 = 9'h49 == first_io_index ? io_grid_73 : _GEN_72; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_74 = 9'h4a == first_io_index ? io_grid_74 : _GEN_73; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_75 = 9'h4b == first_io_index ? io_grid_75 : _GEN_74; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_76 = 9'h4c == first_io_index ? io_grid_76 : _GEN_75; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_77 = 9'h4d == first_io_index ? io_grid_77 : _GEN_76; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_78 = 9'h4e == first_io_index ? io_grid_78 : _GEN_77; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_79 = 9'h4f == first_io_index ? io_grid_79 : _GEN_78; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_80 = 9'h50 == first_io_index ? io_grid_80 : _GEN_79; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_81 = 9'h51 == first_io_index ? io_grid_81 : _GEN_80; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_82 = 9'h52 == first_io_index ? io_grid_82 : _GEN_81; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_83 = 9'h53 == first_io_index ? io_grid_83 : _GEN_82; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_84 = 9'h54 == first_io_index ? io_grid_84 : _GEN_83; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_85 = 9'h55 == first_io_index ? io_grid_85 : _GEN_84; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_86 = 9'h56 == first_io_index ? io_grid_86 : _GEN_85; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_87 = 9'h57 == first_io_index ? io_grid_87 : _GEN_86; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_88 = 9'h58 == first_io_index ? io_grid_88 : _GEN_87; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_89 = 9'h59 == first_io_index ? io_grid_89 : _GEN_88; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_90 = 9'h5a == first_io_index ? io_grid_90 : _GEN_89; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_91 = 9'h5b == first_io_index ? io_grid_91 : _GEN_90; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_92 = 9'h5c == first_io_index ? io_grid_92 : _GEN_91; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_93 = 9'h5d == first_io_index ? io_grid_93 : _GEN_92; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_94 = 9'h5e == first_io_index ? io_grid_94 : _GEN_93; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_95 = 9'h5f == first_io_index ? io_grid_95 : _GEN_94; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_96 = 9'h60 == first_io_index ? io_grid_96 : _GEN_95; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_97 = 9'h61 == first_io_index ? io_grid_97 : _GEN_96; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_98 = 9'h62 == first_io_index ? io_grid_98 : _GEN_97; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_99 = 9'h63 == first_io_index ? io_grid_99 : _GEN_98; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_100 = 9'h64 == first_io_index ? io_grid_100 : _GEN_99; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_101 = 9'h65 == first_io_index ? io_grid_101 : _GEN_100; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_102 = 9'h66 == first_io_index ? io_grid_102 : _GEN_101; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_103 = 9'h67 == first_io_index ? io_grid_103 : _GEN_102; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_104 = 9'h68 == first_io_index ? io_grid_104 : _GEN_103; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_105 = 9'h69 == first_io_index ? io_grid_105 : _GEN_104; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_106 = 9'h6a == first_io_index ? io_grid_106 : _GEN_105; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_107 = 9'h6b == first_io_index ? io_grid_107 : _GEN_106; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_108 = 9'h6c == first_io_index ? io_grid_108 : _GEN_107; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_109 = 9'h6d == first_io_index ? io_grid_109 : _GEN_108; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_110 = 9'h6e == first_io_index ? io_grid_110 : _GEN_109; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_111 = 9'h6f == first_io_index ? io_grid_111 : _GEN_110; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_112 = 9'h70 == first_io_index ? io_grid_112 : _GEN_111; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_113 = 9'h71 == first_io_index ? io_grid_113 : _GEN_112; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_114 = 9'h72 == first_io_index ? io_grid_114 : _GEN_113; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_115 = 9'h73 == first_io_index ? io_grid_115 : _GEN_114; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_116 = 9'h74 == first_io_index ? io_grid_116 : _GEN_115; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_117 = 9'h75 == first_io_index ? io_grid_117 : _GEN_116; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_118 = 9'h76 == first_io_index ? io_grid_118 : _GEN_117; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_119 = 9'h77 == first_io_index ? io_grid_119 : _GEN_118; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_120 = 9'h78 == first_io_index ? io_grid_120 : _GEN_119; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_121 = 9'h79 == first_io_index ? io_grid_121 : _GEN_120; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_122 = 9'h7a == first_io_index ? io_grid_122 : _GEN_121; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_123 = 9'h7b == first_io_index ? io_grid_123 : _GEN_122; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_124 = 9'h7c == first_io_index ? io_grid_124 : _GEN_123; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_125 = 9'h7d == first_io_index ? io_grid_125 : _GEN_124; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_126 = 9'h7e == first_io_index ? io_grid_126 : _GEN_125; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_127 = 9'h7f == first_io_index ? io_grid_127 : _GEN_126; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_128 = 9'h80 == first_io_index ? io_grid_128 : _GEN_127; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_129 = 9'h81 == first_io_index ? io_grid_129 : _GEN_128; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_130 = 9'h82 == first_io_index ? io_grid_130 : _GEN_129; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_131 = 9'h83 == first_io_index ? io_grid_131 : _GEN_130; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_132 = 9'h84 == first_io_index ? io_grid_132 : _GEN_131; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_133 = 9'h85 == first_io_index ? io_grid_133 : _GEN_132; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_134 = 9'h86 == first_io_index ? io_grid_134 : _GEN_133; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_135 = 9'h87 == first_io_index ? io_grid_135 : _GEN_134; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_136 = 9'h88 == first_io_index ? io_grid_136 : _GEN_135; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_137 = 9'h89 == first_io_index ? io_grid_137 : _GEN_136; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_138 = 9'h8a == first_io_index ? io_grid_138 : _GEN_137; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_139 = 9'h8b == first_io_index ? io_grid_139 : _GEN_138; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_140 = 9'h8c == first_io_index ? io_grid_140 : _GEN_139; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_141 = 9'h8d == first_io_index ? io_grid_141 : _GEN_140; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_142 = 9'h8e == first_io_index ? io_grid_142 : _GEN_141; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_143 = 9'h8f == first_io_index ? io_grid_143 : _GEN_142; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_144 = 9'h90 == first_io_index ? io_grid_144 : _GEN_143; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_145 = 9'h91 == first_io_index ? io_grid_145 : _GEN_144; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_146 = 9'h92 == first_io_index ? io_grid_146 : _GEN_145; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_147 = 9'h93 == first_io_index ? io_grid_147 : _GEN_146; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_148 = 9'h94 == first_io_index ? io_grid_148 : _GEN_147; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_149 = 9'h95 == first_io_index ? io_grid_149 : _GEN_148; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_150 = 9'h96 == first_io_index ? io_grid_150 : _GEN_149; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_151 = 9'h97 == first_io_index ? io_grid_151 : _GEN_150; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_152 = 9'h98 == first_io_index ? io_grid_152 : _GEN_151; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_153 = 9'h99 == first_io_index ? io_grid_153 : _GEN_152; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_154 = 9'h9a == first_io_index ? io_grid_154 : _GEN_153; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_155 = 9'h9b == first_io_index ? io_grid_155 : _GEN_154; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_156 = 9'h9c == first_io_index ? io_grid_156 : _GEN_155; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_157 = 9'h9d == first_io_index ? io_grid_157 : _GEN_156; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_158 = 9'h9e == first_io_index ? io_grid_158 : _GEN_157; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_159 = 9'h9f == first_io_index ? io_grid_159 : _GEN_158; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_160 = 9'ha0 == first_io_index ? io_grid_160 : _GEN_159; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_161 = 9'ha1 == first_io_index ? io_grid_161 : _GEN_160; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_162 = 9'ha2 == first_io_index ? io_grid_162 : _GEN_161; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_163 = 9'ha3 == first_io_index ? io_grid_163 : _GEN_162; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_164 = 9'ha4 == first_io_index ? io_grid_164 : _GEN_163; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_165 = 9'ha5 == first_io_index ? io_grid_165 : _GEN_164; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_166 = 9'ha6 == first_io_index ? io_grid_166 : _GEN_165; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_167 = 9'ha7 == first_io_index ? io_grid_167 : _GEN_166; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_168 = 9'ha8 == first_io_index ? io_grid_168 : _GEN_167; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_169 = 9'ha9 == first_io_index ? io_grid_169 : _GEN_168; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_170 = 9'haa == first_io_index ? io_grid_170 : _GEN_169; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_171 = 9'hab == first_io_index ? io_grid_171 : _GEN_170; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_172 = 9'hac == first_io_index ? io_grid_172 : _GEN_171; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_173 = 9'had == first_io_index ? io_grid_173 : _GEN_172; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_174 = 9'hae == first_io_index ? io_grid_174 : _GEN_173; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_175 = 9'haf == first_io_index ? io_grid_175 : _GEN_174; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_176 = 9'hb0 == first_io_index ? io_grid_176 : _GEN_175; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_177 = 9'hb1 == first_io_index ? io_grid_177 : _GEN_176; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_178 = 9'hb2 == first_io_index ? io_grid_178 : _GEN_177; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_179 = 9'hb3 == first_io_index ? io_grid_179 : _GEN_178; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_180 = 9'hb4 == first_io_index ? io_grid_180 : _GEN_179; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_181 = 9'hb5 == first_io_index ? io_grid_181 : _GEN_180; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_182 = 9'hb6 == first_io_index ? io_grid_182 : _GEN_181; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_183 = 9'hb7 == first_io_index ? io_grid_183 : _GEN_182; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_184 = 9'hb8 == first_io_index ? io_grid_184 : _GEN_183; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_185 = 9'hb9 == first_io_index ? io_grid_185 : _GEN_184; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_186 = 9'hba == first_io_index ? io_grid_186 : _GEN_185; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_187 = 9'hbb == first_io_index ? io_grid_187 : _GEN_186; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_188 = 9'hbc == first_io_index ? io_grid_188 : _GEN_187; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_189 = 9'hbd == first_io_index ? io_grid_189 : _GEN_188; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_190 = 9'hbe == first_io_index ? io_grid_190 : _GEN_189; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_191 = 9'hbf == first_io_index ? io_grid_191 : _GEN_190; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_192 = 9'hc0 == first_io_index ? io_grid_192 : _GEN_191; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_193 = 9'hc1 == first_io_index ? io_grid_193 : _GEN_192; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_194 = 9'hc2 == first_io_index ? io_grid_194 : _GEN_193; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_195 = 9'hc3 == first_io_index ? io_grid_195 : _GEN_194; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_196 = 9'hc4 == first_io_index ? io_grid_196 : _GEN_195; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_197 = 9'hc5 == first_io_index ? io_grid_197 : _GEN_196; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_198 = 9'hc6 == first_io_index ? io_grid_198 : _GEN_197; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_199 = 9'hc7 == first_io_index ? io_grid_199 : _GEN_198; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_200 = 9'hc8 == first_io_index ? io_grid_200 : _GEN_199; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_201 = 9'hc9 == first_io_index ? io_grid_201 : _GEN_200; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_202 = 9'hca == first_io_index ? io_grid_202 : _GEN_201; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_203 = 9'hcb == first_io_index ? io_grid_203 : _GEN_202; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_204 = 9'hcc == first_io_index ? io_grid_204 : _GEN_203; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_205 = 9'hcd == first_io_index ? io_grid_205 : _GEN_204; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_206 = 9'hce == first_io_index ? io_grid_206 : _GEN_205; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_207 = 9'hcf == first_io_index ? io_grid_207 : _GEN_206; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_208 = 9'hd0 == first_io_index ? io_grid_208 : _GEN_207; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_209 = 9'hd1 == first_io_index ? io_grid_209 : _GEN_208; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_210 = 9'hd2 == first_io_index ? io_grid_210 : _GEN_209; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_211 = 9'hd3 == first_io_index ? io_grid_211 : _GEN_210; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_212 = 9'hd4 == first_io_index ? io_grid_212 : _GEN_211; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_213 = 9'hd5 == first_io_index ? io_grid_213 : _GEN_212; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_214 = 9'hd6 == first_io_index ? io_grid_214 : _GEN_213; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_215 = 9'hd7 == first_io_index ? io_grid_215 : _GEN_214; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_216 = 9'hd8 == first_io_index ? io_grid_216 : _GEN_215; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_217 = 9'hd9 == first_io_index ? io_grid_217 : _GEN_216; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_218 = 9'hda == first_io_index ? io_grid_218 : _GEN_217; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_219 = 9'hdb == first_io_index ? io_grid_219 : _GEN_218; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_220 = 9'hdc == first_io_index ? io_grid_220 : _GEN_219; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_221 = 9'hdd == first_io_index ? io_grid_221 : _GEN_220; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_222 = 9'hde == first_io_index ? io_grid_222 : _GEN_221; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_223 = 9'hdf == first_io_index ? io_grid_223 : _GEN_222; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_224 = 9'he0 == first_io_index ? io_grid_224 : _GEN_223; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_225 = 9'he1 == first_io_index ? io_grid_225 : _GEN_224; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_226 = 9'he2 == first_io_index ? io_grid_226 : _GEN_225; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_227 = 9'he3 == first_io_index ? io_grid_227 : _GEN_226; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_228 = 9'he4 == first_io_index ? io_grid_228 : _GEN_227; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_229 = 9'he5 == first_io_index ? io_grid_229 : _GEN_228; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_230 = 9'he6 == first_io_index ? io_grid_230 : _GEN_229; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_231 = 9'he7 == first_io_index ? io_grid_231 : _GEN_230; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_232 = 9'he8 == first_io_index ? io_grid_232 : _GEN_231; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_233 = 9'he9 == first_io_index ? io_grid_233 : _GEN_232; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_234 = 9'hea == first_io_index ? io_grid_234 : _GEN_233; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_235 = 9'heb == first_io_index ? io_grid_235 : _GEN_234; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_236 = 9'hec == first_io_index ? io_grid_236 : _GEN_235; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_237 = 9'hed == first_io_index ? io_grid_237 : _GEN_236; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_238 = 9'hee == first_io_index ? io_grid_238 : _GEN_237; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_239 = 9'hef == first_io_index ? io_grid_239 : _GEN_238; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_240 = 9'hf0 == first_io_index ? io_grid_240 : _GEN_239; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_241 = 9'hf1 == first_io_index ? io_grid_241 : _GEN_240; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_242 = 9'hf2 == first_io_index ? io_grid_242 : _GEN_241; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_243 = 9'hf3 == first_io_index ? io_grid_243 : _GEN_242; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_244 = 9'hf4 == first_io_index ? io_grid_244 : _GEN_243; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_245 = 9'hf5 == first_io_index ? io_grid_245 : _GEN_244; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_246 = 9'hf6 == first_io_index ? io_grid_246 : _GEN_245; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_247 = 9'hf7 == first_io_index ? io_grid_247 : _GEN_246; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_248 = 9'hf8 == first_io_index ? io_grid_248 : _GEN_247; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_249 = 9'hf9 == first_io_index ? io_grid_249 : _GEN_248; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_250 = 9'hfa == first_io_index ? io_grid_250 : _GEN_249; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_251 = 9'hfb == first_io_index ? io_grid_251 : _GEN_250; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_252 = 9'hfc == first_io_index ? io_grid_252 : _GEN_251; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_253 = 9'hfd == first_io_index ? io_grid_253 : _GEN_252; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_254 = 9'hfe == first_io_index ? io_grid_254 : _GEN_253; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_255 = 9'hff == first_io_index ? io_grid_255 : _GEN_254; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_256 = 9'h100 == first_io_index ? io_grid_256 : _GEN_255; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_257 = 9'h101 == first_io_index ? io_grid_257 : _GEN_256; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_258 = 9'h102 == first_io_index ? io_grid_258 : _GEN_257; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_259 = 9'h103 == first_io_index ? io_grid_259 : _GEN_258; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_260 = 9'h104 == first_io_index ? io_grid_260 : _GEN_259; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_261 = 9'h105 == first_io_index ? io_grid_261 : _GEN_260; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_262 = 9'h106 == first_io_index ? io_grid_262 : _GEN_261; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_263 = 9'h107 == first_io_index ? io_grid_263 : _GEN_262; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_264 = 9'h108 == first_io_index ? io_grid_264 : _GEN_263; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_265 = 9'h109 == first_io_index ? io_grid_265 : _GEN_264; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_266 = 9'h10a == first_io_index ? io_grid_266 : _GEN_265; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_267 = 9'h10b == first_io_index ? io_grid_267 : _GEN_266; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_268 = 9'h10c == first_io_index ? io_grid_268 : _GEN_267; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_269 = 9'h10d == first_io_index ? io_grid_269 : _GEN_268; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_270 = 9'h10e == first_io_index ? io_grid_270 : _GEN_269; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_271 = 9'h10f == first_io_index ? io_grid_271 : _GEN_270; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_272 = 9'h110 == first_io_index ? io_grid_272 : _GEN_271; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_273 = 9'h111 == first_io_index ? io_grid_273 : _GEN_272; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_274 = 9'h112 == first_io_index ? io_grid_274 : _GEN_273; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_275 = 9'h113 == first_io_index ? io_grid_275 : _GEN_274; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_276 = 9'h114 == first_io_index ? io_grid_276 : _GEN_275; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_277 = 9'h115 == first_io_index ? io_grid_277 : _GEN_276; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_278 = 9'h116 == first_io_index ? io_grid_278 : _GEN_277; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_279 = 9'h117 == first_io_index ? io_grid_279 : _GEN_278; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_280 = 9'h118 == first_io_index ? io_grid_280 : _GEN_279; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_281 = 9'h119 == first_io_index ? io_grid_281 : _GEN_280; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_282 = 9'h11a == first_io_index ? io_grid_282 : _GEN_281; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_283 = 9'h11b == first_io_index ? io_grid_283 : _GEN_282; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_284 = 9'h11c == first_io_index ? io_grid_284 : _GEN_283; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_285 = 9'h11d == first_io_index ? io_grid_285 : _GEN_284; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_286 = 9'h11e == first_io_index ? io_grid_286 : _GEN_285; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_287 = 9'h11f == first_io_index ? io_grid_287 : _GEN_286; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_288 = 9'h120 == first_io_index ? io_grid_288 : _GEN_287; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_289 = 9'h121 == first_io_index ? io_grid_289 : _GEN_288; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_290 = 9'h122 == first_io_index ? io_grid_290 : _GEN_289; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_291 = 9'h123 == first_io_index ? io_grid_291 : _GEN_290; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_292 = 9'h124 == first_io_index ? io_grid_292 : _GEN_291; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_293 = 9'h125 == first_io_index ? io_grid_293 : _GEN_292; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_294 = 9'h126 == first_io_index ? io_grid_294 : _GEN_293; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_295 = 9'h127 == first_io_index ? io_grid_295 : _GEN_294; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_296 = 9'h128 == first_io_index ? io_grid_296 : _GEN_295; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_297 = 9'h129 == first_io_index ? io_grid_297 : _GEN_296; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_298 = 9'h12a == first_io_index ? io_grid_298 : _GEN_297; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire [2:0] _GEN_299 = 9'h12b == first_io_index ? io_grid_299 : _GEN_298; // @[\\src\\main\\scala\\CollisionDetector.scala 34:{50,50}]
  wire  firstCollision = ~(_GEN_299 == 3'h0); // @[\\src\\main\\scala\\CollisionDetector.scala 34:24]
  wire [2:0] _GEN_301 = 9'h1 == second_io_index ? io_grid_1 : io_grid_0; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_302 = 9'h2 == second_io_index ? io_grid_2 : _GEN_301; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_303 = 9'h3 == second_io_index ? io_grid_3 : _GEN_302; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_304 = 9'h4 == second_io_index ? io_grid_4 : _GEN_303; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_305 = 9'h5 == second_io_index ? io_grid_5 : _GEN_304; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_306 = 9'h6 == second_io_index ? io_grid_6 : _GEN_305; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_307 = 9'h7 == second_io_index ? io_grid_7 : _GEN_306; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_308 = 9'h8 == second_io_index ? io_grid_8 : _GEN_307; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_309 = 9'h9 == second_io_index ? io_grid_9 : _GEN_308; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_310 = 9'ha == second_io_index ? io_grid_10 : _GEN_309; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_311 = 9'hb == second_io_index ? io_grid_11 : _GEN_310; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_312 = 9'hc == second_io_index ? io_grid_12 : _GEN_311; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_313 = 9'hd == second_io_index ? io_grid_13 : _GEN_312; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_314 = 9'he == second_io_index ? io_grid_14 : _GEN_313; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_315 = 9'hf == second_io_index ? io_grid_15 : _GEN_314; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_316 = 9'h10 == second_io_index ? io_grid_16 : _GEN_315; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_317 = 9'h11 == second_io_index ? io_grid_17 : _GEN_316; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_318 = 9'h12 == second_io_index ? io_grid_18 : _GEN_317; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_319 = 9'h13 == second_io_index ? io_grid_19 : _GEN_318; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_320 = 9'h14 == second_io_index ? io_grid_20 : _GEN_319; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_321 = 9'h15 == second_io_index ? io_grid_21 : _GEN_320; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_322 = 9'h16 == second_io_index ? io_grid_22 : _GEN_321; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_323 = 9'h17 == second_io_index ? io_grid_23 : _GEN_322; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_324 = 9'h18 == second_io_index ? io_grid_24 : _GEN_323; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_325 = 9'h19 == second_io_index ? io_grid_25 : _GEN_324; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_326 = 9'h1a == second_io_index ? io_grid_26 : _GEN_325; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_327 = 9'h1b == second_io_index ? io_grid_27 : _GEN_326; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_328 = 9'h1c == second_io_index ? io_grid_28 : _GEN_327; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_329 = 9'h1d == second_io_index ? io_grid_29 : _GEN_328; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_330 = 9'h1e == second_io_index ? io_grid_30 : _GEN_329; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_331 = 9'h1f == second_io_index ? io_grid_31 : _GEN_330; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_332 = 9'h20 == second_io_index ? io_grid_32 : _GEN_331; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_333 = 9'h21 == second_io_index ? io_grid_33 : _GEN_332; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_334 = 9'h22 == second_io_index ? io_grid_34 : _GEN_333; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_335 = 9'h23 == second_io_index ? io_grid_35 : _GEN_334; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_336 = 9'h24 == second_io_index ? io_grid_36 : _GEN_335; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_337 = 9'h25 == second_io_index ? io_grid_37 : _GEN_336; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_338 = 9'h26 == second_io_index ? io_grid_38 : _GEN_337; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_339 = 9'h27 == second_io_index ? io_grid_39 : _GEN_338; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_340 = 9'h28 == second_io_index ? io_grid_40 : _GEN_339; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_341 = 9'h29 == second_io_index ? io_grid_41 : _GEN_340; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_342 = 9'h2a == second_io_index ? io_grid_42 : _GEN_341; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_343 = 9'h2b == second_io_index ? io_grid_43 : _GEN_342; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_344 = 9'h2c == second_io_index ? io_grid_44 : _GEN_343; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_345 = 9'h2d == second_io_index ? io_grid_45 : _GEN_344; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_346 = 9'h2e == second_io_index ? io_grid_46 : _GEN_345; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_347 = 9'h2f == second_io_index ? io_grid_47 : _GEN_346; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_348 = 9'h30 == second_io_index ? io_grid_48 : _GEN_347; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_349 = 9'h31 == second_io_index ? io_grid_49 : _GEN_348; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_350 = 9'h32 == second_io_index ? io_grid_50 : _GEN_349; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_351 = 9'h33 == second_io_index ? io_grid_51 : _GEN_350; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_352 = 9'h34 == second_io_index ? io_grid_52 : _GEN_351; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_353 = 9'h35 == second_io_index ? io_grid_53 : _GEN_352; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_354 = 9'h36 == second_io_index ? io_grid_54 : _GEN_353; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_355 = 9'h37 == second_io_index ? io_grid_55 : _GEN_354; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_356 = 9'h38 == second_io_index ? io_grid_56 : _GEN_355; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_357 = 9'h39 == second_io_index ? io_grid_57 : _GEN_356; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_358 = 9'h3a == second_io_index ? io_grid_58 : _GEN_357; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_359 = 9'h3b == second_io_index ? io_grid_59 : _GEN_358; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_360 = 9'h3c == second_io_index ? io_grid_60 : _GEN_359; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_361 = 9'h3d == second_io_index ? io_grid_61 : _GEN_360; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_362 = 9'h3e == second_io_index ? io_grid_62 : _GEN_361; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_363 = 9'h3f == second_io_index ? io_grid_63 : _GEN_362; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_364 = 9'h40 == second_io_index ? io_grid_64 : _GEN_363; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_365 = 9'h41 == second_io_index ? io_grid_65 : _GEN_364; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_366 = 9'h42 == second_io_index ? io_grid_66 : _GEN_365; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_367 = 9'h43 == second_io_index ? io_grid_67 : _GEN_366; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_368 = 9'h44 == second_io_index ? io_grid_68 : _GEN_367; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_369 = 9'h45 == second_io_index ? io_grid_69 : _GEN_368; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_370 = 9'h46 == second_io_index ? io_grid_70 : _GEN_369; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_371 = 9'h47 == second_io_index ? io_grid_71 : _GEN_370; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_372 = 9'h48 == second_io_index ? io_grid_72 : _GEN_371; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_373 = 9'h49 == second_io_index ? io_grid_73 : _GEN_372; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_374 = 9'h4a == second_io_index ? io_grid_74 : _GEN_373; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_375 = 9'h4b == second_io_index ? io_grid_75 : _GEN_374; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_376 = 9'h4c == second_io_index ? io_grid_76 : _GEN_375; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_377 = 9'h4d == second_io_index ? io_grid_77 : _GEN_376; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_378 = 9'h4e == second_io_index ? io_grid_78 : _GEN_377; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_379 = 9'h4f == second_io_index ? io_grid_79 : _GEN_378; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_380 = 9'h50 == second_io_index ? io_grid_80 : _GEN_379; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_381 = 9'h51 == second_io_index ? io_grid_81 : _GEN_380; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_382 = 9'h52 == second_io_index ? io_grid_82 : _GEN_381; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_383 = 9'h53 == second_io_index ? io_grid_83 : _GEN_382; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_384 = 9'h54 == second_io_index ? io_grid_84 : _GEN_383; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_385 = 9'h55 == second_io_index ? io_grid_85 : _GEN_384; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_386 = 9'h56 == second_io_index ? io_grid_86 : _GEN_385; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_387 = 9'h57 == second_io_index ? io_grid_87 : _GEN_386; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_388 = 9'h58 == second_io_index ? io_grid_88 : _GEN_387; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_389 = 9'h59 == second_io_index ? io_grid_89 : _GEN_388; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_390 = 9'h5a == second_io_index ? io_grid_90 : _GEN_389; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_391 = 9'h5b == second_io_index ? io_grid_91 : _GEN_390; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_392 = 9'h5c == second_io_index ? io_grid_92 : _GEN_391; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_393 = 9'h5d == second_io_index ? io_grid_93 : _GEN_392; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_394 = 9'h5e == second_io_index ? io_grid_94 : _GEN_393; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_395 = 9'h5f == second_io_index ? io_grid_95 : _GEN_394; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_396 = 9'h60 == second_io_index ? io_grid_96 : _GEN_395; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_397 = 9'h61 == second_io_index ? io_grid_97 : _GEN_396; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_398 = 9'h62 == second_io_index ? io_grid_98 : _GEN_397; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_399 = 9'h63 == second_io_index ? io_grid_99 : _GEN_398; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_400 = 9'h64 == second_io_index ? io_grid_100 : _GEN_399; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_401 = 9'h65 == second_io_index ? io_grid_101 : _GEN_400; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_402 = 9'h66 == second_io_index ? io_grid_102 : _GEN_401; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_403 = 9'h67 == second_io_index ? io_grid_103 : _GEN_402; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_404 = 9'h68 == second_io_index ? io_grid_104 : _GEN_403; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_405 = 9'h69 == second_io_index ? io_grid_105 : _GEN_404; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_406 = 9'h6a == second_io_index ? io_grid_106 : _GEN_405; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_407 = 9'h6b == second_io_index ? io_grid_107 : _GEN_406; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_408 = 9'h6c == second_io_index ? io_grid_108 : _GEN_407; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_409 = 9'h6d == second_io_index ? io_grid_109 : _GEN_408; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_410 = 9'h6e == second_io_index ? io_grid_110 : _GEN_409; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_411 = 9'h6f == second_io_index ? io_grid_111 : _GEN_410; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_412 = 9'h70 == second_io_index ? io_grid_112 : _GEN_411; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_413 = 9'h71 == second_io_index ? io_grid_113 : _GEN_412; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_414 = 9'h72 == second_io_index ? io_grid_114 : _GEN_413; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_415 = 9'h73 == second_io_index ? io_grid_115 : _GEN_414; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_416 = 9'h74 == second_io_index ? io_grid_116 : _GEN_415; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_417 = 9'h75 == second_io_index ? io_grid_117 : _GEN_416; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_418 = 9'h76 == second_io_index ? io_grid_118 : _GEN_417; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_419 = 9'h77 == second_io_index ? io_grid_119 : _GEN_418; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_420 = 9'h78 == second_io_index ? io_grid_120 : _GEN_419; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_421 = 9'h79 == second_io_index ? io_grid_121 : _GEN_420; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_422 = 9'h7a == second_io_index ? io_grid_122 : _GEN_421; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_423 = 9'h7b == second_io_index ? io_grid_123 : _GEN_422; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_424 = 9'h7c == second_io_index ? io_grid_124 : _GEN_423; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_425 = 9'h7d == second_io_index ? io_grid_125 : _GEN_424; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_426 = 9'h7e == second_io_index ? io_grid_126 : _GEN_425; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_427 = 9'h7f == second_io_index ? io_grid_127 : _GEN_426; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_428 = 9'h80 == second_io_index ? io_grid_128 : _GEN_427; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_429 = 9'h81 == second_io_index ? io_grid_129 : _GEN_428; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_430 = 9'h82 == second_io_index ? io_grid_130 : _GEN_429; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_431 = 9'h83 == second_io_index ? io_grid_131 : _GEN_430; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_432 = 9'h84 == second_io_index ? io_grid_132 : _GEN_431; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_433 = 9'h85 == second_io_index ? io_grid_133 : _GEN_432; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_434 = 9'h86 == second_io_index ? io_grid_134 : _GEN_433; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_435 = 9'h87 == second_io_index ? io_grid_135 : _GEN_434; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_436 = 9'h88 == second_io_index ? io_grid_136 : _GEN_435; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_437 = 9'h89 == second_io_index ? io_grid_137 : _GEN_436; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_438 = 9'h8a == second_io_index ? io_grid_138 : _GEN_437; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_439 = 9'h8b == second_io_index ? io_grid_139 : _GEN_438; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_440 = 9'h8c == second_io_index ? io_grid_140 : _GEN_439; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_441 = 9'h8d == second_io_index ? io_grid_141 : _GEN_440; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_442 = 9'h8e == second_io_index ? io_grid_142 : _GEN_441; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_443 = 9'h8f == second_io_index ? io_grid_143 : _GEN_442; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_444 = 9'h90 == second_io_index ? io_grid_144 : _GEN_443; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_445 = 9'h91 == second_io_index ? io_grid_145 : _GEN_444; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_446 = 9'h92 == second_io_index ? io_grid_146 : _GEN_445; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_447 = 9'h93 == second_io_index ? io_grid_147 : _GEN_446; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_448 = 9'h94 == second_io_index ? io_grid_148 : _GEN_447; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_449 = 9'h95 == second_io_index ? io_grid_149 : _GEN_448; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_450 = 9'h96 == second_io_index ? io_grid_150 : _GEN_449; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_451 = 9'h97 == second_io_index ? io_grid_151 : _GEN_450; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_452 = 9'h98 == second_io_index ? io_grid_152 : _GEN_451; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_453 = 9'h99 == second_io_index ? io_grid_153 : _GEN_452; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_454 = 9'h9a == second_io_index ? io_grid_154 : _GEN_453; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_455 = 9'h9b == second_io_index ? io_grid_155 : _GEN_454; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_456 = 9'h9c == second_io_index ? io_grid_156 : _GEN_455; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_457 = 9'h9d == second_io_index ? io_grid_157 : _GEN_456; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_458 = 9'h9e == second_io_index ? io_grid_158 : _GEN_457; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_459 = 9'h9f == second_io_index ? io_grid_159 : _GEN_458; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_460 = 9'ha0 == second_io_index ? io_grid_160 : _GEN_459; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_461 = 9'ha1 == second_io_index ? io_grid_161 : _GEN_460; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_462 = 9'ha2 == second_io_index ? io_grid_162 : _GEN_461; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_463 = 9'ha3 == second_io_index ? io_grid_163 : _GEN_462; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_464 = 9'ha4 == second_io_index ? io_grid_164 : _GEN_463; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_465 = 9'ha5 == second_io_index ? io_grid_165 : _GEN_464; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_466 = 9'ha6 == second_io_index ? io_grid_166 : _GEN_465; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_467 = 9'ha7 == second_io_index ? io_grid_167 : _GEN_466; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_468 = 9'ha8 == second_io_index ? io_grid_168 : _GEN_467; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_469 = 9'ha9 == second_io_index ? io_grid_169 : _GEN_468; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_470 = 9'haa == second_io_index ? io_grid_170 : _GEN_469; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_471 = 9'hab == second_io_index ? io_grid_171 : _GEN_470; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_472 = 9'hac == second_io_index ? io_grid_172 : _GEN_471; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_473 = 9'had == second_io_index ? io_grid_173 : _GEN_472; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_474 = 9'hae == second_io_index ? io_grid_174 : _GEN_473; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_475 = 9'haf == second_io_index ? io_grid_175 : _GEN_474; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_476 = 9'hb0 == second_io_index ? io_grid_176 : _GEN_475; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_477 = 9'hb1 == second_io_index ? io_grid_177 : _GEN_476; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_478 = 9'hb2 == second_io_index ? io_grid_178 : _GEN_477; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_479 = 9'hb3 == second_io_index ? io_grid_179 : _GEN_478; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_480 = 9'hb4 == second_io_index ? io_grid_180 : _GEN_479; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_481 = 9'hb5 == second_io_index ? io_grid_181 : _GEN_480; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_482 = 9'hb6 == second_io_index ? io_grid_182 : _GEN_481; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_483 = 9'hb7 == second_io_index ? io_grid_183 : _GEN_482; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_484 = 9'hb8 == second_io_index ? io_grid_184 : _GEN_483; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_485 = 9'hb9 == second_io_index ? io_grid_185 : _GEN_484; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_486 = 9'hba == second_io_index ? io_grid_186 : _GEN_485; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_487 = 9'hbb == second_io_index ? io_grid_187 : _GEN_486; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_488 = 9'hbc == second_io_index ? io_grid_188 : _GEN_487; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_489 = 9'hbd == second_io_index ? io_grid_189 : _GEN_488; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_490 = 9'hbe == second_io_index ? io_grid_190 : _GEN_489; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_491 = 9'hbf == second_io_index ? io_grid_191 : _GEN_490; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_492 = 9'hc0 == second_io_index ? io_grid_192 : _GEN_491; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_493 = 9'hc1 == second_io_index ? io_grid_193 : _GEN_492; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_494 = 9'hc2 == second_io_index ? io_grid_194 : _GEN_493; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_495 = 9'hc3 == second_io_index ? io_grid_195 : _GEN_494; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_496 = 9'hc4 == second_io_index ? io_grid_196 : _GEN_495; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_497 = 9'hc5 == second_io_index ? io_grid_197 : _GEN_496; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_498 = 9'hc6 == second_io_index ? io_grid_198 : _GEN_497; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_499 = 9'hc7 == second_io_index ? io_grid_199 : _GEN_498; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_500 = 9'hc8 == second_io_index ? io_grid_200 : _GEN_499; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_501 = 9'hc9 == second_io_index ? io_grid_201 : _GEN_500; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_502 = 9'hca == second_io_index ? io_grid_202 : _GEN_501; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_503 = 9'hcb == second_io_index ? io_grid_203 : _GEN_502; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_504 = 9'hcc == second_io_index ? io_grid_204 : _GEN_503; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_505 = 9'hcd == second_io_index ? io_grid_205 : _GEN_504; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_506 = 9'hce == second_io_index ? io_grid_206 : _GEN_505; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_507 = 9'hcf == second_io_index ? io_grid_207 : _GEN_506; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_508 = 9'hd0 == second_io_index ? io_grid_208 : _GEN_507; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_509 = 9'hd1 == second_io_index ? io_grid_209 : _GEN_508; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_510 = 9'hd2 == second_io_index ? io_grid_210 : _GEN_509; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_511 = 9'hd3 == second_io_index ? io_grid_211 : _GEN_510; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_512 = 9'hd4 == second_io_index ? io_grid_212 : _GEN_511; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_513 = 9'hd5 == second_io_index ? io_grid_213 : _GEN_512; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_514 = 9'hd6 == second_io_index ? io_grid_214 : _GEN_513; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_515 = 9'hd7 == second_io_index ? io_grid_215 : _GEN_514; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_516 = 9'hd8 == second_io_index ? io_grid_216 : _GEN_515; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_517 = 9'hd9 == second_io_index ? io_grid_217 : _GEN_516; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_518 = 9'hda == second_io_index ? io_grid_218 : _GEN_517; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_519 = 9'hdb == second_io_index ? io_grid_219 : _GEN_518; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_520 = 9'hdc == second_io_index ? io_grid_220 : _GEN_519; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_521 = 9'hdd == second_io_index ? io_grid_221 : _GEN_520; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_522 = 9'hde == second_io_index ? io_grid_222 : _GEN_521; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_523 = 9'hdf == second_io_index ? io_grid_223 : _GEN_522; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_524 = 9'he0 == second_io_index ? io_grid_224 : _GEN_523; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_525 = 9'he1 == second_io_index ? io_grid_225 : _GEN_524; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_526 = 9'he2 == second_io_index ? io_grid_226 : _GEN_525; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_527 = 9'he3 == second_io_index ? io_grid_227 : _GEN_526; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_528 = 9'he4 == second_io_index ? io_grid_228 : _GEN_527; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_529 = 9'he5 == second_io_index ? io_grid_229 : _GEN_528; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_530 = 9'he6 == second_io_index ? io_grid_230 : _GEN_529; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_531 = 9'he7 == second_io_index ? io_grid_231 : _GEN_530; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_532 = 9'he8 == second_io_index ? io_grid_232 : _GEN_531; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_533 = 9'he9 == second_io_index ? io_grid_233 : _GEN_532; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_534 = 9'hea == second_io_index ? io_grid_234 : _GEN_533; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_535 = 9'heb == second_io_index ? io_grid_235 : _GEN_534; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_536 = 9'hec == second_io_index ? io_grid_236 : _GEN_535; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_537 = 9'hed == second_io_index ? io_grid_237 : _GEN_536; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_538 = 9'hee == second_io_index ? io_grid_238 : _GEN_537; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_539 = 9'hef == second_io_index ? io_grid_239 : _GEN_538; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_540 = 9'hf0 == second_io_index ? io_grid_240 : _GEN_539; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_541 = 9'hf1 == second_io_index ? io_grid_241 : _GEN_540; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_542 = 9'hf2 == second_io_index ? io_grid_242 : _GEN_541; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_543 = 9'hf3 == second_io_index ? io_grid_243 : _GEN_542; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_544 = 9'hf4 == second_io_index ? io_grid_244 : _GEN_543; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_545 = 9'hf5 == second_io_index ? io_grid_245 : _GEN_544; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_546 = 9'hf6 == second_io_index ? io_grid_246 : _GEN_545; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_547 = 9'hf7 == second_io_index ? io_grid_247 : _GEN_546; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_548 = 9'hf8 == second_io_index ? io_grid_248 : _GEN_547; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_549 = 9'hf9 == second_io_index ? io_grid_249 : _GEN_548; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_550 = 9'hfa == second_io_index ? io_grid_250 : _GEN_549; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_551 = 9'hfb == second_io_index ? io_grid_251 : _GEN_550; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_552 = 9'hfc == second_io_index ? io_grid_252 : _GEN_551; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_553 = 9'hfd == second_io_index ? io_grid_253 : _GEN_552; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_554 = 9'hfe == second_io_index ? io_grid_254 : _GEN_553; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_555 = 9'hff == second_io_index ? io_grid_255 : _GEN_554; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_556 = 9'h100 == second_io_index ? io_grid_256 : _GEN_555; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_557 = 9'h101 == second_io_index ? io_grid_257 : _GEN_556; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_558 = 9'h102 == second_io_index ? io_grid_258 : _GEN_557; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_559 = 9'h103 == second_io_index ? io_grid_259 : _GEN_558; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_560 = 9'h104 == second_io_index ? io_grid_260 : _GEN_559; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_561 = 9'h105 == second_io_index ? io_grid_261 : _GEN_560; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_562 = 9'h106 == second_io_index ? io_grid_262 : _GEN_561; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_563 = 9'h107 == second_io_index ? io_grid_263 : _GEN_562; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_564 = 9'h108 == second_io_index ? io_grid_264 : _GEN_563; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_565 = 9'h109 == second_io_index ? io_grid_265 : _GEN_564; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_566 = 9'h10a == second_io_index ? io_grid_266 : _GEN_565; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_567 = 9'h10b == second_io_index ? io_grid_267 : _GEN_566; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_568 = 9'h10c == second_io_index ? io_grid_268 : _GEN_567; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_569 = 9'h10d == second_io_index ? io_grid_269 : _GEN_568; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_570 = 9'h10e == second_io_index ? io_grid_270 : _GEN_569; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_571 = 9'h10f == second_io_index ? io_grid_271 : _GEN_570; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_572 = 9'h110 == second_io_index ? io_grid_272 : _GEN_571; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_573 = 9'h111 == second_io_index ? io_grid_273 : _GEN_572; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_574 = 9'h112 == second_io_index ? io_grid_274 : _GEN_573; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_575 = 9'h113 == second_io_index ? io_grid_275 : _GEN_574; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_576 = 9'h114 == second_io_index ? io_grid_276 : _GEN_575; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_577 = 9'h115 == second_io_index ? io_grid_277 : _GEN_576; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_578 = 9'h116 == second_io_index ? io_grid_278 : _GEN_577; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_579 = 9'h117 == second_io_index ? io_grid_279 : _GEN_578; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_580 = 9'h118 == second_io_index ? io_grid_280 : _GEN_579; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_581 = 9'h119 == second_io_index ? io_grid_281 : _GEN_580; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_582 = 9'h11a == second_io_index ? io_grid_282 : _GEN_581; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_583 = 9'h11b == second_io_index ? io_grid_283 : _GEN_582; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_584 = 9'h11c == second_io_index ? io_grid_284 : _GEN_583; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_585 = 9'h11d == second_io_index ? io_grid_285 : _GEN_584; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_586 = 9'h11e == second_io_index ? io_grid_286 : _GEN_585; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_587 = 9'h11f == second_io_index ? io_grid_287 : _GEN_586; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_588 = 9'h120 == second_io_index ? io_grid_288 : _GEN_587; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_589 = 9'h121 == second_io_index ? io_grid_289 : _GEN_588; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_590 = 9'h122 == second_io_index ? io_grid_290 : _GEN_589; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_591 = 9'h123 == second_io_index ? io_grid_291 : _GEN_590; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_592 = 9'h124 == second_io_index ? io_grid_292 : _GEN_591; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_593 = 9'h125 == second_io_index ? io_grid_293 : _GEN_592; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_594 = 9'h126 == second_io_index ? io_grid_294 : _GEN_593; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_595 = 9'h127 == second_io_index ? io_grid_295 : _GEN_594; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_596 = 9'h128 == second_io_index ? io_grid_296 : _GEN_595; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_597 = 9'h129 == second_io_index ? io_grid_297 : _GEN_596; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_598 = 9'h12a == second_io_index ? io_grid_298 : _GEN_597; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire [2:0] _GEN_599 = 9'h12b == second_io_index ? io_grid_299 : _GEN_598; // @[\\src\\main\\scala\\CollisionDetector.scala 35:{52,52}]
  wire  secondCollision = ~(_GEN_599 == 3'h0); // @[\\src\\main\\scala\\CollisionDetector.scala 35:25]
  wire [2:0] _GEN_601 = 9'h1 == third_io_index ? io_grid_1 : io_grid_0; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_602 = 9'h2 == third_io_index ? io_grid_2 : _GEN_601; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_603 = 9'h3 == third_io_index ? io_grid_3 : _GEN_602; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_604 = 9'h4 == third_io_index ? io_grid_4 : _GEN_603; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_605 = 9'h5 == third_io_index ? io_grid_5 : _GEN_604; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_606 = 9'h6 == third_io_index ? io_grid_6 : _GEN_605; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_607 = 9'h7 == third_io_index ? io_grid_7 : _GEN_606; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_608 = 9'h8 == third_io_index ? io_grid_8 : _GEN_607; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_609 = 9'h9 == third_io_index ? io_grid_9 : _GEN_608; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_610 = 9'ha == third_io_index ? io_grid_10 : _GEN_609; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_611 = 9'hb == third_io_index ? io_grid_11 : _GEN_610; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_612 = 9'hc == third_io_index ? io_grid_12 : _GEN_611; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_613 = 9'hd == third_io_index ? io_grid_13 : _GEN_612; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_614 = 9'he == third_io_index ? io_grid_14 : _GEN_613; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_615 = 9'hf == third_io_index ? io_grid_15 : _GEN_614; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_616 = 9'h10 == third_io_index ? io_grid_16 : _GEN_615; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_617 = 9'h11 == third_io_index ? io_grid_17 : _GEN_616; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_618 = 9'h12 == third_io_index ? io_grid_18 : _GEN_617; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_619 = 9'h13 == third_io_index ? io_grid_19 : _GEN_618; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_620 = 9'h14 == third_io_index ? io_grid_20 : _GEN_619; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_621 = 9'h15 == third_io_index ? io_grid_21 : _GEN_620; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_622 = 9'h16 == third_io_index ? io_grid_22 : _GEN_621; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_623 = 9'h17 == third_io_index ? io_grid_23 : _GEN_622; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_624 = 9'h18 == third_io_index ? io_grid_24 : _GEN_623; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_625 = 9'h19 == third_io_index ? io_grid_25 : _GEN_624; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_626 = 9'h1a == third_io_index ? io_grid_26 : _GEN_625; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_627 = 9'h1b == third_io_index ? io_grid_27 : _GEN_626; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_628 = 9'h1c == third_io_index ? io_grid_28 : _GEN_627; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_629 = 9'h1d == third_io_index ? io_grid_29 : _GEN_628; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_630 = 9'h1e == third_io_index ? io_grid_30 : _GEN_629; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_631 = 9'h1f == third_io_index ? io_grid_31 : _GEN_630; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_632 = 9'h20 == third_io_index ? io_grid_32 : _GEN_631; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_633 = 9'h21 == third_io_index ? io_grid_33 : _GEN_632; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_634 = 9'h22 == third_io_index ? io_grid_34 : _GEN_633; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_635 = 9'h23 == third_io_index ? io_grid_35 : _GEN_634; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_636 = 9'h24 == third_io_index ? io_grid_36 : _GEN_635; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_637 = 9'h25 == third_io_index ? io_grid_37 : _GEN_636; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_638 = 9'h26 == third_io_index ? io_grid_38 : _GEN_637; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_639 = 9'h27 == third_io_index ? io_grid_39 : _GEN_638; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_640 = 9'h28 == third_io_index ? io_grid_40 : _GEN_639; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_641 = 9'h29 == third_io_index ? io_grid_41 : _GEN_640; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_642 = 9'h2a == third_io_index ? io_grid_42 : _GEN_641; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_643 = 9'h2b == third_io_index ? io_grid_43 : _GEN_642; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_644 = 9'h2c == third_io_index ? io_grid_44 : _GEN_643; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_645 = 9'h2d == third_io_index ? io_grid_45 : _GEN_644; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_646 = 9'h2e == third_io_index ? io_grid_46 : _GEN_645; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_647 = 9'h2f == third_io_index ? io_grid_47 : _GEN_646; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_648 = 9'h30 == third_io_index ? io_grid_48 : _GEN_647; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_649 = 9'h31 == third_io_index ? io_grid_49 : _GEN_648; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_650 = 9'h32 == third_io_index ? io_grid_50 : _GEN_649; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_651 = 9'h33 == third_io_index ? io_grid_51 : _GEN_650; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_652 = 9'h34 == third_io_index ? io_grid_52 : _GEN_651; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_653 = 9'h35 == third_io_index ? io_grid_53 : _GEN_652; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_654 = 9'h36 == third_io_index ? io_grid_54 : _GEN_653; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_655 = 9'h37 == third_io_index ? io_grid_55 : _GEN_654; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_656 = 9'h38 == third_io_index ? io_grid_56 : _GEN_655; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_657 = 9'h39 == third_io_index ? io_grid_57 : _GEN_656; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_658 = 9'h3a == third_io_index ? io_grid_58 : _GEN_657; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_659 = 9'h3b == third_io_index ? io_grid_59 : _GEN_658; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_660 = 9'h3c == third_io_index ? io_grid_60 : _GEN_659; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_661 = 9'h3d == third_io_index ? io_grid_61 : _GEN_660; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_662 = 9'h3e == third_io_index ? io_grid_62 : _GEN_661; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_663 = 9'h3f == third_io_index ? io_grid_63 : _GEN_662; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_664 = 9'h40 == third_io_index ? io_grid_64 : _GEN_663; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_665 = 9'h41 == third_io_index ? io_grid_65 : _GEN_664; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_666 = 9'h42 == third_io_index ? io_grid_66 : _GEN_665; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_667 = 9'h43 == third_io_index ? io_grid_67 : _GEN_666; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_668 = 9'h44 == third_io_index ? io_grid_68 : _GEN_667; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_669 = 9'h45 == third_io_index ? io_grid_69 : _GEN_668; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_670 = 9'h46 == third_io_index ? io_grid_70 : _GEN_669; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_671 = 9'h47 == third_io_index ? io_grid_71 : _GEN_670; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_672 = 9'h48 == third_io_index ? io_grid_72 : _GEN_671; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_673 = 9'h49 == third_io_index ? io_grid_73 : _GEN_672; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_674 = 9'h4a == third_io_index ? io_grid_74 : _GEN_673; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_675 = 9'h4b == third_io_index ? io_grid_75 : _GEN_674; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_676 = 9'h4c == third_io_index ? io_grid_76 : _GEN_675; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_677 = 9'h4d == third_io_index ? io_grid_77 : _GEN_676; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_678 = 9'h4e == third_io_index ? io_grid_78 : _GEN_677; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_679 = 9'h4f == third_io_index ? io_grid_79 : _GEN_678; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_680 = 9'h50 == third_io_index ? io_grid_80 : _GEN_679; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_681 = 9'h51 == third_io_index ? io_grid_81 : _GEN_680; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_682 = 9'h52 == third_io_index ? io_grid_82 : _GEN_681; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_683 = 9'h53 == third_io_index ? io_grid_83 : _GEN_682; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_684 = 9'h54 == third_io_index ? io_grid_84 : _GEN_683; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_685 = 9'h55 == third_io_index ? io_grid_85 : _GEN_684; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_686 = 9'h56 == third_io_index ? io_grid_86 : _GEN_685; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_687 = 9'h57 == third_io_index ? io_grid_87 : _GEN_686; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_688 = 9'h58 == third_io_index ? io_grid_88 : _GEN_687; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_689 = 9'h59 == third_io_index ? io_grid_89 : _GEN_688; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_690 = 9'h5a == third_io_index ? io_grid_90 : _GEN_689; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_691 = 9'h5b == third_io_index ? io_grid_91 : _GEN_690; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_692 = 9'h5c == third_io_index ? io_grid_92 : _GEN_691; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_693 = 9'h5d == third_io_index ? io_grid_93 : _GEN_692; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_694 = 9'h5e == third_io_index ? io_grid_94 : _GEN_693; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_695 = 9'h5f == third_io_index ? io_grid_95 : _GEN_694; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_696 = 9'h60 == third_io_index ? io_grid_96 : _GEN_695; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_697 = 9'h61 == third_io_index ? io_grid_97 : _GEN_696; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_698 = 9'h62 == third_io_index ? io_grid_98 : _GEN_697; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_699 = 9'h63 == third_io_index ? io_grid_99 : _GEN_698; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_700 = 9'h64 == third_io_index ? io_grid_100 : _GEN_699; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_701 = 9'h65 == third_io_index ? io_grid_101 : _GEN_700; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_702 = 9'h66 == third_io_index ? io_grid_102 : _GEN_701; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_703 = 9'h67 == third_io_index ? io_grid_103 : _GEN_702; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_704 = 9'h68 == third_io_index ? io_grid_104 : _GEN_703; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_705 = 9'h69 == third_io_index ? io_grid_105 : _GEN_704; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_706 = 9'h6a == third_io_index ? io_grid_106 : _GEN_705; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_707 = 9'h6b == third_io_index ? io_grid_107 : _GEN_706; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_708 = 9'h6c == third_io_index ? io_grid_108 : _GEN_707; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_709 = 9'h6d == third_io_index ? io_grid_109 : _GEN_708; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_710 = 9'h6e == third_io_index ? io_grid_110 : _GEN_709; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_711 = 9'h6f == third_io_index ? io_grid_111 : _GEN_710; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_712 = 9'h70 == third_io_index ? io_grid_112 : _GEN_711; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_713 = 9'h71 == third_io_index ? io_grid_113 : _GEN_712; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_714 = 9'h72 == third_io_index ? io_grid_114 : _GEN_713; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_715 = 9'h73 == third_io_index ? io_grid_115 : _GEN_714; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_716 = 9'h74 == third_io_index ? io_grid_116 : _GEN_715; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_717 = 9'h75 == third_io_index ? io_grid_117 : _GEN_716; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_718 = 9'h76 == third_io_index ? io_grid_118 : _GEN_717; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_719 = 9'h77 == third_io_index ? io_grid_119 : _GEN_718; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_720 = 9'h78 == third_io_index ? io_grid_120 : _GEN_719; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_721 = 9'h79 == third_io_index ? io_grid_121 : _GEN_720; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_722 = 9'h7a == third_io_index ? io_grid_122 : _GEN_721; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_723 = 9'h7b == third_io_index ? io_grid_123 : _GEN_722; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_724 = 9'h7c == third_io_index ? io_grid_124 : _GEN_723; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_725 = 9'h7d == third_io_index ? io_grid_125 : _GEN_724; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_726 = 9'h7e == third_io_index ? io_grid_126 : _GEN_725; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_727 = 9'h7f == third_io_index ? io_grid_127 : _GEN_726; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_728 = 9'h80 == third_io_index ? io_grid_128 : _GEN_727; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_729 = 9'h81 == third_io_index ? io_grid_129 : _GEN_728; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_730 = 9'h82 == third_io_index ? io_grid_130 : _GEN_729; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_731 = 9'h83 == third_io_index ? io_grid_131 : _GEN_730; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_732 = 9'h84 == third_io_index ? io_grid_132 : _GEN_731; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_733 = 9'h85 == third_io_index ? io_grid_133 : _GEN_732; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_734 = 9'h86 == third_io_index ? io_grid_134 : _GEN_733; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_735 = 9'h87 == third_io_index ? io_grid_135 : _GEN_734; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_736 = 9'h88 == third_io_index ? io_grid_136 : _GEN_735; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_737 = 9'h89 == third_io_index ? io_grid_137 : _GEN_736; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_738 = 9'h8a == third_io_index ? io_grid_138 : _GEN_737; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_739 = 9'h8b == third_io_index ? io_grid_139 : _GEN_738; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_740 = 9'h8c == third_io_index ? io_grid_140 : _GEN_739; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_741 = 9'h8d == third_io_index ? io_grid_141 : _GEN_740; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_742 = 9'h8e == third_io_index ? io_grid_142 : _GEN_741; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_743 = 9'h8f == third_io_index ? io_grid_143 : _GEN_742; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_744 = 9'h90 == third_io_index ? io_grid_144 : _GEN_743; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_745 = 9'h91 == third_io_index ? io_grid_145 : _GEN_744; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_746 = 9'h92 == third_io_index ? io_grid_146 : _GEN_745; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_747 = 9'h93 == third_io_index ? io_grid_147 : _GEN_746; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_748 = 9'h94 == third_io_index ? io_grid_148 : _GEN_747; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_749 = 9'h95 == third_io_index ? io_grid_149 : _GEN_748; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_750 = 9'h96 == third_io_index ? io_grid_150 : _GEN_749; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_751 = 9'h97 == third_io_index ? io_grid_151 : _GEN_750; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_752 = 9'h98 == third_io_index ? io_grid_152 : _GEN_751; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_753 = 9'h99 == third_io_index ? io_grid_153 : _GEN_752; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_754 = 9'h9a == third_io_index ? io_grid_154 : _GEN_753; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_755 = 9'h9b == third_io_index ? io_grid_155 : _GEN_754; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_756 = 9'h9c == third_io_index ? io_grid_156 : _GEN_755; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_757 = 9'h9d == third_io_index ? io_grid_157 : _GEN_756; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_758 = 9'h9e == third_io_index ? io_grid_158 : _GEN_757; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_759 = 9'h9f == third_io_index ? io_grid_159 : _GEN_758; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_760 = 9'ha0 == third_io_index ? io_grid_160 : _GEN_759; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_761 = 9'ha1 == third_io_index ? io_grid_161 : _GEN_760; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_762 = 9'ha2 == third_io_index ? io_grid_162 : _GEN_761; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_763 = 9'ha3 == third_io_index ? io_grid_163 : _GEN_762; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_764 = 9'ha4 == third_io_index ? io_grid_164 : _GEN_763; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_765 = 9'ha5 == third_io_index ? io_grid_165 : _GEN_764; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_766 = 9'ha6 == third_io_index ? io_grid_166 : _GEN_765; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_767 = 9'ha7 == third_io_index ? io_grid_167 : _GEN_766; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_768 = 9'ha8 == third_io_index ? io_grid_168 : _GEN_767; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_769 = 9'ha9 == third_io_index ? io_grid_169 : _GEN_768; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_770 = 9'haa == third_io_index ? io_grid_170 : _GEN_769; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_771 = 9'hab == third_io_index ? io_grid_171 : _GEN_770; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_772 = 9'hac == third_io_index ? io_grid_172 : _GEN_771; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_773 = 9'had == third_io_index ? io_grid_173 : _GEN_772; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_774 = 9'hae == third_io_index ? io_grid_174 : _GEN_773; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_775 = 9'haf == third_io_index ? io_grid_175 : _GEN_774; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_776 = 9'hb0 == third_io_index ? io_grid_176 : _GEN_775; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_777 = 9'hb1 == third_io_index ? io_grid_177 : _GEN_776; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_778 = 9'hb2 == third_io_index ? io_grid_178 : _GEN_777; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_779 = 9'hb3 == third_io_index ? io_grid_179 : _GEN_778; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_780 = 9'hb4 == third_io_index ? io_grid_180 : _GEN_779; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_781 = 9'hb5 == third_io_index ? io_grid_181 : _GEN_780; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_782 = 9'hb6 == third_io_index ? io_grid_182 : _GEN_781; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_783 = 9'hb7 == third_io_index ? io_grid_183 : _GEN_782; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_784 = 9'hb8 == third_io_index ? io_grid_184 : _GEN_783; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_785 = 9'hb9 == third_io_index ? io_grid_185 : _GEN_784; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_786 = 9'hba == third_io_index ? io_grid_186 : _GEN_785; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_787 = 9'hbb == third_io_index ? io_grid_187 : _GEN_786; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_788 = 9'hbc == third_io_index ? io_grid_188 : _GEN_787; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_789 = 9'hbd == third_io_index ? io_grid_189 : _GEN_788; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_790 = 9'hbe == third_io_index ? io_grid_190 : _GEN_789; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_791 = 9'hbf == third_io_index ? io_grid_191 : _GEN_790; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_792 = 9'hc0 == third_io_index ? io_grid_192 : _GEN_791; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_793 = 9'hc1 == third_io_index ? io_grid_193 : _GEN_792; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_794 = 9'hc2 == third_io_index ? io_grid_194 : _GEN_793; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_795 = 9'hc3 == third_io_index ? io_grid_195 : _GEN_794; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_796 = 9'hc4 == third_io_index ? io_grid_196 : _GEN_795; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_797 = 9'hc5 == third_io_index ? io_grid_197 : _GEN_796; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_798 = 9'hc6 == third_io_index ? io_grid_198 : _GEN_797; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_799 = 9'hc7 == third_io_index ? io_grid_199 : _GEN_798; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_800 = 9'hc8 == third_io_index ? io_grid_200 : _GEN_799; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_801 = 9'hc9 == third_io_index ? io_grid_201 : _GEN_800; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_802 = 9'hca == third_io_index ? io_grid_202 : _GEN_801; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_803 = 9'hcb == third_io_index ? io_grid_203 : _GEN_802; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_804 = 9'hcc == third_io_index ? io_grid_204 : _GEN_803; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_805 = 9'hcd == third_io_index ? io_grid_205 : _GEN_804; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_806 = 9'hce == third_io_index ? io_grid_206 : _GEN_805; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_807 = 9'hcf == third_io_index ? io_grid_207 : _GEN_806; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_808 = 9'hd0 == third_io_index ? io_grid_208 : _GEN_807; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_809 = 9'hd1 == third_io_index ? io_grid_209 : _GEN_808; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_810 = 9'hd2 == third_io_index ? io_grid_210 : _GEN_809; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_811 = 9'hd3 == third_io_index ? io_grid_211 : _GEN_810; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_812 = 9'hd4 == third_io_index ? io_grid_212 : _GEN_811; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_813 = 9'hd5 == third_io_index ? io_grid_213 : _GEN_812; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_814 = 9'hd6 == third_io_index ? io_grid_214 : _GEN_813; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_815 = 9'hd7 == third_io_index ? io_grid_215 : _GEN_814; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_816 = 9'hd8 == third_io_index ? io_grid_216 : _GEN_815; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_817 = 9'hd9 == third_io_index ? io_grid_217 : _GEN_816; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_818 = 9'hda == third_io_index ? io_grid_218 : _GEN_817; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_819 = 9'hdb == third_io_index ? io_grid_219 : _GEN_818; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_820 = 9'hdc == third_io_index ? io_grid_220 : _GEN_819; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_821 = 9'hdd == third_io_index ? io_grid_221 : _GEN_820; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_822 = 9'hde == third_io_index ? io_grid_222 : _GEN_821; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_823 = 9'hdf == third_io_index ? io_grid_223 : _GEN_822; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_824 = 9'he0 == third_io_index ? io_grid_224 : _GEN_823; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_825 = 9'he1 == third_io_index ? io_grid_225 : _GEN_824; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_826 = 9'he2 == third_io_index ? io_grid_226 : _GEN_825; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_827 = 9'he3 == third_io_index ? io_grid_227 : _GEN_826; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_828 = 9'he4 == third_io_index ? io_grid_228 : _GEN_827; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_829 = 9'he5 == third_io_index ? io_grid_229 : _GEN_828; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_830 = 9'he6 == third_io_index ? io_grid_230 : _GEN_829; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_831 = 9'he7 == third_io_index ? io_grid_231 : _GEN_830; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_832 = 9'he8 == third_io_index ? io_grid_232 : _GEN_831; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_833 = 9'he9 == third_io_index ? io_grid_233 : _GEN_832; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_834 = 9'hea == third_io_index ? io_grid_234 : _GEN_833; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_835 = 9'heb == third_io_index ? io_grid_235 : _GEN_834; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_836 = 9'hec == third_io_index ? io_grid_236 : _GEN_835; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_837 = 9'hed == third_io_index ? io_grid_237 : _GEN_836; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_838 = 9'hee == third_io_index ? io_grid_238 : _GEN_837; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_839 = 9'hef == third_io_index ? io_grid_239 : _GEN_838; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_840 = 9'hf0 == third_io_index ? io_grid_240 : _GEN_839; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_841 = 9'hf1 == third_io_index ? io_grid_241 : _GEN_840; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_842 = 9'hf2 == third_io_index ? io_grid_242 : _GEN_841; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_843 = 9'hf3 == third_io_index ? io_grid_243 : _GEN_842; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_844 = 9'hf4 == third_io_index ? io_grid_244 : _GEN_843; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_845 = 9'hf5 == third_io_index ? io_grid_245 : _GEN_844; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_846 = 9'hf6 == third_io_index ? io_grid_246 : _GEN_845; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_847 = 9'hf7 == third_io_index ? io_grid_247 : _GEN_846; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_848 = 9'hf8 == third_io_index ? io_grid_248 : _GEN_847; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_849 = 9'hf9 == third_io_index ? io_grid_249 : _GEN_848; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_850 = 9'hfa == third_io_index ? io_grid_250 : _GEN_849; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_851 = 9'hfb == third_io_index ? io_grid_251 : _GEN_850; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_852 = 9'hfc == third_io_index ? io_grid_252 : _GEN_851; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_853 = 9'hfd == third_io_index ? io_grid_253 : _GEN_852; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_854 = 9'hfe == third_io_index ? io_grid_254 : _GEN_853; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_855 = 9'hff == third_io_index ? io_grid_255 : _GEN_854; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_856 = 9'h100 == third_io_index ? io_grid_256 : _GEN_855; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_857 = 9'h101 == third_io_index ? io_grid_257 : _GEN_856; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_858 = 9'h102 == third_io_index ? io_grid_258 : _GEN_857; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_859 = 9'h103 == third_io_index ? io_grid_259 : _GEN_858; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_860 = 9'h104 == third_io_index ? io_grid_260 : _GEN_859; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_861 = 9'h105 == third_io_index ? io_grid_261 : _GEN_860; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_862 = 9'h106 == third_io_index ? io_grid_262 : _GEN_861; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_863 = 9'h107 == third_io_index ? io_grid_263 : _GEN_862; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_864 = 9'h108 == third_io_index ? io_grid_264 : _GEN_863; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_865 = 9'h109 == third_io_index ? io_grid_265 : _GEN_864; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_866 = 9'h10a == third_io_index ? io_grid_266 : _GEN_865; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_867 = 9'h10b == third_io_index ? io_grid_267 : _GEN_866; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_868 = 9'h10c == third_io_index ? io_grid_268 : _GEN_867; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_869 = 9'h10d == third_io_index ? io_grid_269 : _GEN_868; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_870 = 9'h10e == third_io_index ? io_grid_270 : _GEN_869; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_871 = 9'h10f == third_io_index ? io_grid_271 : _GEN_870; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_872 = 9'h110 == third_io_index ? io_grid_272 : _GEN_871; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_873 = 9'h111 == third_io_index ? io_grid_273 : _GEN_872; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_874 = 9'h112 == third_io_index ? io_grid_274 : _GEN_873; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_875 = 9'h113 == third_io_index ? io_grid_275 : _GEN_874; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_876 = 9'h114 == third_io_index ? io_grid_276 : _GEN_875; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_877 = 9'h115 == third_io_index ? io_grid_277 : _GEN_876; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_878 = 9'h116 == third_io_index ? io_grid_278 : _GEN_877; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_879 = 9'h117 == third_io_index ? io_grid_279 : _GEN_878; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_880 = 9'h118 == third_io_index ? io_grid_280 : _GEN_879; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_881 = 9'h119 == third_io_index ? io_grid_281 : _GEN_880; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_882 = 9'h11a == third_io_index ? io_grid_282 : _GEN_881; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_883 = 9'h11b == third_io_index ? io_grid_283 : _GEN_882; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_884 = 9'h11c == third_io_index ? io_grid_284 : _GEN_883; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_885 = 9'h11d == third_io_index ? io_grid_285 : _GEN_884; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_886 = 9'h11e == third_io_index ? io_grid_286 : _GEN_885; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_887 = 9'h11f == third_io_index ? io_grid_287 : _GEN_886; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_888 = 9'h120 == third_io_index ? io_grid_288 : _GEN_887; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_889 = 9'h121 == third_io_index ? io_grid_289 : _GEN_888; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_890 = 9'h122 == third_io_index ? io_grid_290 : _GEN_889; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_891 = 9'h123 == third_io_index ? io_grid_291 : _GEN_890; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_892 = 9'h124 == third_io_index ? io_grid_292 : _GEN_891; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_893 = 9'h125 == third_io_index ? io_grid_293 : _GEN_892; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_894 = 9'h126 == third_io_index ? io_grid_294 : _GEN_893; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_895 = 9'h127 == third_io_index ? io_grid_295 : _GEN_894; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_896 = 9'h128 == third_io_index ? io_grid_296 : _GEN_895; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_897 = 9'h129 == third_io_index ? io_grid_297 : _GEN_896; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_898 = 9'h12a == third_io_index ? io_grid_298 : _GEN_897; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire [2:0] _GEN_899 = 9'h12b == third_io_index ? io_grid_299 : _GEN_898; // @[\\src\\main\\scala\\CollisionDetector.scala 36:{50,50}]
  wire  thirdCollision = ~(_GEN_899 == 3'h0); // @[\\src\\main\\scala\\CollisionDetector.scala 36:24]
  wire [2:0] _GEN_901 = 9'h1 == fourth_io_index ? io_grid_1 : io_grid_0; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_902 = 9'h2 == fourth_io_index ? io_grid_2 : _GEN_901; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_903 = 9'h3 == fourth_io_index ? io_grid_3 : _GEN_902; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_904 = 9'h4 == fourth_io_index ? io_grid_4 : _GEN_903; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_905 = 9'h5 == fourth_io_index ? io_grid_5 : _GEN_904; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_906 = 9'h6 == fourth_io_index ? io_grid_6 : _GEN_905; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_907 = 9'h7 == fourth_io_index ? io_grid_7 : _GEN_906; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_908 = 9'h8 == fourth_io_index ? io_grid_8 : _GEN_907; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_909 = 9'h9 == fourth_io_index ? io_grid_9 : _GEN_908; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_910 = 9'ha == fourth_io_index ? io_grid_10 : _GEN_909; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_911 = 9'hb == fourth_io_index ? io_grid_11 : _GEN_910; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_912 = 9'hc == fourth_io_index ? io_grid_12 : _GEN_911; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_913 = 9'hd == fourth_io_index ? io_grid_13 : _GEN_912; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_914 = 9'he == fourth_io_index ? io_grid_14 : _GEN_913; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_915 = 9'hf == fourth_io_index ? io_grid_15 : _GEN_914; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_916 = 9'h10 == fourth_io_index ? io_grid_16 : _GEN_915; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_917 = 9'h11 == fourth_io_index ? io_grid_17 : _GEN_916; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_918 = 9'h12 == fourth_io_index ? io_grid_18 : _GEN_917; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_919 = 9'h13 == fourth_io_index ? io_grid_19 : _GEN_918; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_920 = 9'h14 == fourth_io_index ? io_grid_20 : _GEN_919; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_921 = 9'h15 == fourth_io_index ? io_grid_21 : _GEN_920; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_922 = 9'h16 == fourth_io_index ? io_grid_22 : _GEN_921; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_923 = 9'h17 == fourth_io_index ? io_grid_23 : _GEN_922; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_924 = 9'h18 == fourth_io_index ? io_grid_24 : _GEN_923; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_925 = 9'h19 == fourth_io_index ? io_grid_25 : _GEN_924; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_926 = 9'h1a == fourth_io_index ? io_grid_26 : _GEN_925; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_927 = 9'h1b == fourth_io_index ? io_grid_27 : _GEN_926; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_928 = 9'h1c == fourth_io_index ? io_grid_28 : _GEN_927; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_929 = 9'h1d == fourth_io_index ? io_grid_29 : _GEN_928; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_930 = 9'h1e == fourth_io_index ? io_grid_30 : _GEN_929; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_931 = 9'h1f == fourth_io_index ? io_grid_31 : _GEN_930; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_932 = 9'h20 == fourth_io_index ? io_grid_32 : _GEN_931; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_933 = 9'h21 == fourth_io_index ? io_grid_33 : _GEN_932; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_934 = 9'h22 == fourth_io_index ? io_grid_34 : _GEN_933; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_935 = 9'h23 == fourth_io_index ? io_grid_35 : _GEN_934; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_936 = 9'h24 == fourth_io_index ? io_grid_36 : _GEN_935; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_937 = 9'h25 == fourth_io_index ? io_grid_37 : _GEN_936; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_938 = 9'h26 == fourth_io_index ? io_grid_38 : _GEN_937; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_939 = 9'h27 == fourth_io_index ? io_grid_39 : _GEN_938; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_940 = 9'h28 == fourth_io_index ? io_grid_40 : _GEN_939; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_941 = 9'h29 == fourth_io_index ? io_grid_41 : _GEN_940; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_942 = 9'h2a == fourth_io_index ? io_grid_42 : _GEN_941; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_943 = 9'h2b == fourth_io_index ? io_grid_43 : _GEN_942; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_944 = 9'h2c == fourth_io_index ? io_grid_44 : _GEN_943; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_945 = 9'h2d == fourth_io_index ? io_grid_45 : _GEN_944; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_946 = 9'h2e == fourth_io_index ? io_grid_46 : _GEN_945; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_947 = 9'h2f == fourth_io_index ? io_grid_47 : _GEN_946; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_948 = 9'h30 == fourth_io_index ? io_grid_48 : _GEN_947; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_949 = 9'h31 == fourth_io_index ? io_grid_49 : _GEN_948; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_950 = 9'h32 == fourth_io_index ? io_grid_50 : _GEN_949; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_951 = 9'h33 == fourth_io_index ? io_grid_51 : _GEN_950; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_952 = 9'h34 == fourth_io_index ? io_grid_52 : _GEN_951; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_953 = 9'h35 == fourth_io_index ? io_grid_53 : _GEN_952; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_954 = 9'h36 == fourth_io_index ? io_grid_54 : _GEN_953; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_955 = 9'h37 == fourth_io_index ? io_grid_55 : _GEN_954; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_956 = 9'h38 == fourth_io_index ? io_grid_56 : _GEN_955; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_957 = 9'h39 == fourth_io_index ? io_grid_57 : _GEN_956; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_958 = 9'h3a == fourth_io_index ? io_grid_58 : _GEN_957; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_959 = 9'h3b == fourth_io_index ? io_grid_59 : _GEN_958; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_960 = 9'h3c == fourth_io_index ? io_grid_60 : _GEN_959; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_961 = 9'h3d == fourth_io_index ? io_grid_61 : _GEN_960; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_962 = 9'h3e == fourth_io_index ? io_grid_62 : _GEN_961; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_963 = 9'h3f == fourth_io_index ? io_grid_63 : _GEN_962; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_964 = 9'h40 == fourth_io_index ? io_grid_64 : _GEN_963; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_965 = 9'h41 == fourth_io_index ? io_grid_65 : _GEN_964; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_966 = 9'h42 == fourth_io_index ? io_grid_66 : _GEN_965; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_967 = 9'h43 == fourth_io_index ? io_grid_67 : _GEN_966; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_968 = 9'h44 == fourth_io_index ? io_grid_68 : _GEN_967; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_969 = 9'h45 == fourth_io_index ? io_grid_69 : _GEN_968; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_970 = 9'h46 == fourth_io_index ? io_grid_70 : _GEN_969; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_971 = 9'h47 == fourth_io_index ? io_grid_71 : _GEN_970; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_972 = 9'h48 == fourth_io_index ? io_grid_72 : _GEN_971; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_973 = 9'h49 == fourth_io_index ? io_grid_73 : _GEN_972; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_974 = 9'h4a == fourth_io_index ? io_grid_74 : _GEN_973; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_975 = 9'h4b == fourth_io_index ? io_grid_75 : _GEN_974; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_976 = 9'h4c == fourth_io_index ? io_grid_76 : _GEN_975; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_977 = 9'h4d == fourth_io_index ? io_grid_77 : _GEN_976; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_978 = 9'h4e == fourth_io_index ? io_grid_78 : _GEN_977; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_979 = 9'h4f == fourth_io_index ? io_grid_79 : _GEN_978; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_980 = 9'h50 == fourth_io_index ? io_grid_80 : _GEN_979; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_981 = 9'h51 == fourth_io_index ? io_grid_81 : _GEN_980; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_982 = 9'h52 == fourth_io_index ? io_grid_82 : _GEN_981; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_983 = 9'h53 == fourth_io_index ? io_grid_83 : _GEN_982; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_984 = 9'h54 == fourth_io_index ? io_grid_84 : _GEN_983; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_985 = 9'h55 == fourth_io_index ? io_grid_85 : _GEN_984; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_986 = 9'h56 == fourth_io_index ? io_grid_86 : _GEN_985; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_987 = 9'h57 == fourth_io_index ? io_grid_87 : _GEN_986; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_988 = 9'h58 == fourth_io_index ? io_grid_88 : _GEN_987; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_989 = 9'h59 == fourth_io_index ? io_grid_89 : _GEN_988; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_990 = 9'h5a == fourth_io_index ? io_grid_90 : _GEN_989; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_991 = 9'h5b == fourth_io_index ? io_grid_91 : _GEN_990; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_992 = 9'h5c == fourth_io_index ? io_grid_92 : _GEN_991; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_993 = 9'h5d == fourth_io_index ? io_grid_93 : _GEN_992; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_994 = 9'h5e == fourth_io_index ? io_grid_94 : _GEN_993; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_995 = 9'h5f == fourth_io_index ? io_grid_95 : _GEN_994; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_996 = 9'h60 == fourth_io_index ? io_grid_96 : _GEN_995; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_997 = 9'h61 == fourth_io_index ? io_grid_97 : _GEN_996; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_998 = 9'h62 == fourth_io_index ? io_grid_98 : _GEN_997; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_999 = 9'h63 == fourth_io_index ? io_grid_99 : _GEN_998; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1000 = 9'h64 == fourth_io_index ? io_grid_100 : _GEN_999; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1001 = 9'h65 == fourth_io_index ? io_grid_101 : _GEN_1000; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1002 = 9'h66 == fourth_io_index ? io_grid_102 : _GEN_1001; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1003 = 9'h67 == fourth_io_index ? io_grid_103 : _GEN_1002; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1004 = 9'h68 == fourth_io_index ? io_grid_104 : _GEN_1003; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1005 = 9'h69 == fourth_io_index ? io_grid_105 : _GEN_1004; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1006 = 9'h6a == fourth_io_index ? io_grid_106 : _GEN_1005; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1007 = 9'h6b == fourth_io_index ? io_grid_107 : _GEN_1006; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1008 = 9'h6c == fourth_io_index ? io_grid_108 : _GEN_1007; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1009 = 9'h6d == fourth_io_index ? io_grid_109 : _GEN_1008; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1010 = 9'h6e == fourth_io_index ? io_grid_110 : _GEN_1009; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1011 = 9'h6f == fourth_io_index ? io_grid_111 : _GEN_1010; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1012 = 9'h70 == fourth_io_index ? io_grid_112 : _GEN_1011; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1013 = 9'h71 == fourth_io_index ? io_grid_113 : _GEN_1012; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1014 = 9'h72 == fourth_io_index ? io_grid_114 : _GEN_1013; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1015 = 9'h73 == fourth_io_index ? io_grid_115 : _GEN_1014; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1016 = 9'h74 == fourth_io_index ? io_grid_116 : _GEN_1015; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1017 = 9'h75 == fourth_io_index ? io_grid_117 : _GEN_1016; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1018 = 9'h76 == fourth_io_index ? io_grid_118 : _GEN_1017; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1019 = 9'h77 == fourth_io_index ? io_grid_119 : _GEN_1018; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1020 = 9'h78 == fourth_io_index ? io_grid_120 : _GEN_1019; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1021 = 9'h79 == fourth_io_index ? io_grid_121 : _GEN_1020; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1022 = 9'h7a == fourth_io_index ? io_grid_122 : _GEN_1021; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1023 = 9'h7b == fourth_io_index ? io_grid_123 : _GEN_1022; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1024 = 9'h7c == fourth_io_index ? io_grid_124 : _GEN_1023; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1025 = 9'h7d == fourth_io_index ? io_grid_125 : _GEN_1024; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1026 = 9'h7e == fourth_io_index ? io_grid_126 : _GEN_1025; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1027 = 9'h7f == fourth_io_index ? io_grid_127 : _GEN_1026; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1028 = 9'h80 == fourth_io_index ? io_grid_128 : _GEN_1027; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1029 = 9'h81 == fourth_io_index ? io_grid_129 : _GEN_1028; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1030 = 9'h82 == fourth_io_index ? io_grid_130 : _GEN_1029; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1031 = 9'h83 == fourth_io_index ? io_grid_131 : _GEN_1030; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1032 = 9'h84 == fourth_io_index ? io_grid_132 : _GEN_1031; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1033 = 9'h85 == fourth_io_index ? io_grid_133 : _GEN_1032; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1034 = 9'h86 == fourth_io_index ? io_grid_134 : _GEN_1033; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1035 = 9'h87 == fourth_io_index ? io_grid_135 : _GEN_1034; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1036 = 9'h88 == fourth_io_index ? io_grid_136 : _GEN_1035; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1037 = 9'h89 == fourth_io_index ? io_grid_137 : _GEN_1036; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1038 = 9'h8a == fourth_io_index ? io_grid_138 : _GEN_1037; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1039 = 9'h8b == fourth_io_index ? io_grid_139 : _GEN_1038; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1040 = 9'h8c == fourth_io_index ? io_grid_140 : _GEN_1039; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1041 = 9'h8d == fourth_io_index ? io_grid_141 : _GEN_1040; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1042 = 9'h8e == fourth_io_index ? io_grid_142 : _GEN_1041; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1043 = 9'h8f == fourth_io_index ? io_grid_143 : _GEN_1042; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1044 = 9'h90 == fourth_io_index ? io_grid_144 : _GEN_1043; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1045 = 9'h91 == fourth_io_index ? io_grid_145 : _GEN_1044; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1046 = 9'h92 == fourth_io_index ? io_grid_146 : _GEN_1045; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1047 = 9'h93 == fourth_io_index ? io_grid_147 : _GEN_1046; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1048 = 9'h94 == fourth_io_index ? io_grid_148 : _GEN_1047; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1049 = 9'h95 == fourth_io_index ? io_grid_149 : _GEN_1048; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1050 = 9'h96 == fourth_io_index ? io_grid_150 : _GEN_1049; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1051 = 9'h97 == fourth_io_index ? io_grid_151 : _GEN_1050; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1052 = 9'h98 == fourth_io_index ? io_grid_152 : _GEN_1051; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1053 = 9'h99 == fourth_io_index ? io_grid_153 : _GEN_1052; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1054 = 9'h9a == fourth_io_index ? io_grid_154 : _GEN_1053; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1055 = 9'h9b == fourth_io_index ? io_grid_155 : _GEN_1054; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1056 = 9'h9c == fourth_io_index ? io_grid_156 : _GEN_1055; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1057 = 9'h9d == fourth_io_index ? io_grid_157 : _GEN_1056; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1058 = 9'h9e == fourth_io_index ? io_grid_158 : _GEN_1057; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1059 = 9'h9f == fourth_io_index ? io_grid_159 : _GEN_1058; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1060 = 9'ha0 == fourth_io_index ? io_grid_160 : _GEN_1059; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1061 = 9'ha1 == fourth_io_index ? io_grid_161 : _GEN_1060; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1062 = 9'ha2 == fourth_io_index ? io_grid_162 : _GEN_1061; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1063 = 9'ha3 == fourth_io_index ? io_grid_163 : _GEN_1062; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1064 = 9'ha4 == fourth_io_index ? io_grid_164 : _GEN_1063; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1065 = 9'ha5 == fourth_io_index ? io_grid_165 : _GEN_1064; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1066 = 9'ha6 == fourth_io_index ? io_grid_166 : _GEN_1065; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1067 = 9'ha7 == fourth_io_index ? io_grid_167 : _GEN_1066; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1068 = 9'ha8 == fourth_io_index ? io_grid_168 : _GEN_1067; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1069 = 9'ha9 == fourth_io_index ? io_grid_169 : _GEN_1068; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1070 = 9'haa == fourth_io_index ? io_grid_170 : _GEN_1069; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1071 = 9'hab == fourth_io_index ? io_grid_171 : _GEN_1070; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1072 = 9'hac == fourth_io_index ? io_grid_172 : _GEN_1071; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1073 = 9'had == fourth_io_index ? io_grid_173 : _GEN_1072; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1074 = 9'hae == fourth_io_index ? io_grid_174 : _GEN_1073; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1075 = 9'haf == fourth_io_index ? io_grid_175 : _GEN_1074; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1076 = 9'hb0 == fourth_io_index ? io_grid_176 : _GEN_1075; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1077 = 9'hb1 == fourth_io_index ? io_grid_177 : _GEN_1076; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1078 = 9'hb2 == fourth_io_index ? io_grid_178 : _GEN_1077; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1079 = 9'hb3 == fourth_io_index ? io_grid_179 : _GEN_1078; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1080 = 9'hb4 == fourth_io_index ? io_grid_180 : _GEN_1079; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1081 = 9'hb5 == fourth_io_index ? io_grid_181 : _GEN_1080; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1082 = 9'hb6 == fourth_io_index ? io_grid_182 : _GEN_1081; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1083 = 9'hb7 == fourth_io_index ? io_grid_183 : _GEN_1082; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1084 = 9'hb8 == fourth_io_index ? io_grid_184 : _GEN_1083; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1085 = 9'hb9 == fourth_io_index ? io_grid_185 : _GEN_1084; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1086 = 9'hba == fourth_io_index ? io_grid_186 : _GEN_1085; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1087 = 9'hbb == fourth_io_index ? io_grid_187 : _GEN_1086; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1088 = 9'hbc == fourth_io_index ? io_grid_188 : _GEN_1087; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1089 = 9'hbd == fourth_io_index ? io_grid_189 : _GEN_1088; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1090 = 9'hbe == fourth_io_index ? io_grid_190 : _GEN_1089; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1091 = 9'hbf == fourth_io_index ? io_grid_191 : _GEN_1090; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1092 = 9'hc0 == fourth_io_index ? io_grid_192 : _GEN_1091; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1093 = 9'hc1 == fourth_io_index ? io_grid_193 : _GEN_1092; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1094 = 9'hc2 == fourth_io_index ? io_grid_194 : _GEN_1093; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1095 = 9'hc3 == fourth_io_index ? io_grid_195 : _GEN_1094; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1096 = 9'hc4 == fourth_io_index ? io_grid_196 : _GEN_1095; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1097 = 9'hc5 == fourth_io_index ? io_grid_197 : _GEN_1096; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1098 = 9'hc6 == fourth_io_index ? io_grid_198 : _GEN_1097; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1099 = 9'hc7 == fourth_io_index ? io_grid_199 : _GEN_1098; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1100 = 9'hc8 == fourth_io_index ? io_grid_200 : _GEN_1099; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1101 = 9'hc9 == fourth_io_index ? io_grid_201 : _GEN_1100; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1102 = 9'hca == fourth_io_index ? io_grid_202 : _GEN_1101; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1103 = 9'hcb == fourth_io_index ? io_grid_203 : _GEN_1102; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1104 = 9'hcc == fourth_io_index ? io_grid_204 : _GEN_1103; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1105 = 9'hcd == fourth_io_index ? io_grid_205 : _GEN_1104; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1106 = 9'hce == fourth_io_index ? io_grid_206 : _GEN_1105; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1107 = 9'hcf == fourth_io_index ? io_grid_207 : _GEN_1106; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1108 = 9'hd0 == fourth_io_index ? io_grid_208 : _GEN_1107; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1109 = 9'hd1 == fourth_io_index ? io_grid_209 : _GEN_1108; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1110 = 9'hd2 == fourth_io_index ? io_grid_210 : _GEN_1109; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1111 = 9'hd3 == fourth_io_index ? io_grid_211 : _GEN_1110; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1112 = 9'hd4 == fourth_io_index ? io_grid_212 : _GEN_1111; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1113 = 9'hd5 == fourth_io_index ? io_grid_213 : _GEN_1112; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1114 = 9'hd6 == fourth_io_index ? io_grid_214 : _GEN_1113; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1115 = 9'hd7 == fourth_io_index ? io_grid_215 : _GEN_1114; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1116 = 9'hd8 == fourth_io_index ? io_grid_216 : _GEN_1115; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1117 = 9'hd9 == fourth_io_index ? io_grid_217 : _GEN_1116; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1118 = 9'hda == fourth_io_index ? io_grid_218 : _GEN_1117; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1119 = 9'hdb == fourth_io_index ? io_grid_219 : _GEN_1118; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1120 = 9'hdc == fourth_io_index ? io_grid_220 : _GEN_1119; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1121 = 9'hdd == fourth_io_index ? io_grid_221 : _GEN_1120; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1122 = 9'hde == fourth_io_index ? io_grid_222 : _GEN_1121; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1123 = 9'hdf == fourth_io_index ? io_grid_223 : _GEN_1122; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1124 = 9'he0 == fourth_io_index ? io_grid_224 : _GEN_1123; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1125 = 9'he1 == fourth_io_index ? io_grid_225 : _GEN_1124; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1126 = 9'he2 == fourth_io_index ? io_grid_226 : _GEN_1125; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1127 = 9'he3 == fourth_io_index ? io_grid_227 : _GEN_1126; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1128 = 9'he4 == fourth_io_index ? io_grid_228 : _GEN_1127; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1129 = 9'he5 == fourth_io_index ? io_grid_229 : _GEN_1128; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1130 = 9'he6 == fourth_io_index ? io_grid_230 : _GEN_1129; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1131 = 9'he7 == fourth_io_index ? io_grid_231 : _GEN_1130; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1132 = 9'he8 == fourth_io_index ? io_grid_232 : _GEN_1131; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1133 = 9'he9 == fourth_io_index ? io_grid_233 : _GEN_1132; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1134 = 9'hea == fourth_io_index ? io_grid_234 : _GEN_1133; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1135 = 9'heb == fourth_io_index ? io_grid_235 : _GEN_1134; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1136 = 9'hec == fourth_io_index ? io_grid_236 : _GEN_1135; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1137 = 9'hed == fourth_io_index ? io_grid_237 : _GEN_1136; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1138 = 9'hee == fourth_io_index ? io_grid_238 : _GEN_1137; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1139 = 9'hef == fourth_io_index ? io_grid_239 : _GEN_1138; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1140 = 9'hf0 == fourth_io_index ? io_grid_240 : _GEN_1139; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1141 = 9'hf1 == fourth_io_index ? io_grid_241 : _GEN_1140; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1142 = 9'hf2 == fourth_io_index ? io_grid_242 : _GEN_1141; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1143 = 9'hf3 == fourth_io_index ? io_grid_243 : _GEN_1142; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1144 = 9'hf4 == fourth_io_index ? io_grid_244 : _GEN_1143; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1145 = 9'hf5 == fourth_io_index ? io_grid_245 : _GEN_1144; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1146 = 9'hf6 == fourth_io_index ? io_grid_246 : _GEN_1145; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1147 = 9'hf7 == fourth_io_index ? io_grid_247 : _GEN_1146; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1148 = 9'hf8 == fourth_io_index ? io_grid_248 : _GEN_1147; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1149 = 9'hf9 == fourth_io_index ? io_grid_249 : _GEN_1148; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1150 = 9'hfa == fourth_io_index ? io_grid_250 : _GEN_1149; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1151 = 9'hfb == fourth_io_index ? io_grid_251 : _GEN_1150; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1152 = 9'hfc == fourth_io_index ? io_grid_252 : _GEN_1151; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1153 = 9'hfd == fourth_io_index ? io_grid_253 : _GEN_1152; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1154 = 9'hfe == fourth_io_index ? io_grid_254 : _GEN_1153; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1155 = 9'hff == fourth_io_index ? io_grid_255 : _GEN_1154; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1156 = 9'h100 == fourth_io_index ? io_grid_256 : _GEN_1155; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1157 = 9'h101 == fourth_io_index ? io_grid_257 : _GEN_1156; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1158 = 9'h102 == fourth_io_index ? io_grid_258 : _GEN_1157; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1159 = 9'h103 == fourth_io_index ? io_grid_259 : _GEN_1158; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1160 = 9'h104 == fourth_io_index ? io_grid_260 : _GEN_1159; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1161 = 9'h105 == fourth_io_index ? io_grid_261 : _GEN_1160; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1162 = 9'h106 == fourth_io_index ? io_grid_262 : _GEN_1161; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1163 = 9'h107 == fourth_io_index ? io_grid_263 : _GEN_1162; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1164 = 9'h108 == fourth_io_index ? io_grid_264 : _GEN_1163; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1165 = 9'h109 == fourth_io_index ? io_grid_265 : _GEN_1164; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1166 = 9'h10a == fourth_io_index ? io_grid_266 : _GEN_1165; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1167 = 9'h10b == fourth_io_index ? io_grid_267 : _GEN_1166; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1168 = 9'h10c == fourth_io_index ? io_grid_268 : _GEN_1167; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1169 = 9'h10d == fourth_io_index ? io_grid_269 : _GEN_1168; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1170 = 9'h10e == fourth_io_index ? io_grid_270 : _GEN_1169; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1171 = 9'h10f == fourth_io_index ? io_grid_271 : _GEN_1170; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1172 = 9'h110 == fourth_io_index ? io_grid_272 : _GEN_1171; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1173 = 9'h111 == fourth_io_index ? io_grid_273 : _GEN_1172; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1174 = 9'h112 == fourth_io_index ? io_grid_274 : _GEN_1173; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1175 = 9'h113 == fourth_io_index ? io_grid_275 : _GEN_1174; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1176 = 9'h114 == fourth_io_index ? io_grid_276 : _GEN_1175; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1177 = 9'h115 == fourth_io_index ? io_grid_277 : _GEN_1176; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1178 = 9'h116 == fourth_io_index ? io_grid_278 : _GEN_1177; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1179 = 9'h117 == fourth_io_index ? io_grid_279 : _GEN_1178; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1180 = 9'h118 == fourth_io_index ? io_grid_280 : _GEN_1179; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1181 = 9'h119 == fourth_io_index ? io_grid_281 : _GEN_1180; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1182 = 9'h11a == fourth_io_index ? io_grid_282 : _GEN_1181; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1183 = 9'h11b == fourth_io_index ? io_grid_283 : _GEN_1182; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1184 = 9'h11c == fourth_io_index ? io_grid_284 : _GEN_1183; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1185 = 9'h11d == fourth_io_index ? io_grid_285 : _GEN_1184; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1186 = 9'h11e == fourth_io_index ? io_grid_286 : _GEN_1185; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1187 = 9'h11f == fourth_io_index ? io_grid_287 : _GEN_1186; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1188 = 9'h120 == fourth_io_index ? io_grid_288 : _GEN_1187; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1189 = 9'h121 == fourth_io_index ? io_grid_289 : _GEN_1188; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1190 = 9'h122 == fourth_io_index ? io_grid_290 : _GEN_1189; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1191 = 9'h123 == fourth_io_index ? io_grid_291 : _GEN_1190; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1192 = 9'h124 == fourth_io_index ? io_grid_292 : _GEN_1191; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1193 = 9'h125 == fourth_io_index ? io_grid_293 : _GEN_1192; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1194 = 9'h126 == fourth_io_index ? io_grid_294 : _GEN_1193; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1195 = 9'h127 == fourth_io_index ? io_grid_295 : _GEN_1194; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1196 = 9'h128 == fourth_io_index ? io_grid_296 : _GEN_1195; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1197 = 9'h129 == fourth_io_index ? io_grid_297 : _GEN_1196; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1198 = 9'h12a == fourth_io_index ? io_grid_298 : _GEN_1197; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire [2:0] _GEN_1199 = 9'h12b == fourth_io_index ? io_grid_299 : _GEN_1198; // @[\\src\\main\\scala\\CollisionDetector.scala 37:{52,52}]
  wire  fourthCollision = ~(_GEN_1199 == 3'h0); // @[\\src\\main\\scala\\CollisionDetector.scala 37:25]
  PosToGridIndex first ( // @[\\src\\main\\scala\\CollisionDetector.scala 22:21]
    .io_xPos(first_io_xPos),
    .io_yPos(first_io_yPos),
    .io_index(first_io_index)
  );
  PosToGridIndex second ( // @[\\src\\main\\scala\\CollisionDetector.scala 23:22]
    .io_xPos(second_io_xPos),
    .io_yPos(second_io_yPos),
    .io_index(second_io_index)
  );
  PosToGridIndex third ( // @[\\src\\main\\scala\\CollisionDetector.scala 24:21]
    .io_xPos(third_io_xPos),
    .io_yPos(third_io_yPos),
    .io_index(third_io_index)
  );
  PosToGridIndex fourth ( // @[\\src\\main\\scala\\CollisionDetector.scala 25:23]
    .io_xPos(fourth_io_xPos),
    .io_yPos(fourth_io_yPos),
    .io_index(fourth_io_index)
  );
  assign io_isCollision = firstCollision | secondCollision | thirdCollision | fourthCollision; // @[\\src\\main\\scala\\CollisionDetector.scala 38:73]
  assign first_io_xPos = $signed(io_xPos) + $signed(_GEN_1200); // @[\\src\\main\\scala\\CollisionDetector.scala 26:28]
  assign first_io_yPos = $signed(io_yPos) + $signed(_GEN_1201); // @[\\src\\main\\scala\\CollisionDetector.scala 27:28]
  assign second_io_xPos = $signed(io_xPos) + $signed(_GEN_1202); // @[\\src\\main\\scala\\CollisionDetector.scala 28:29]
  assign second_io_yPos = $signed(io_yPos) + $signed(_GEN_1203); // @[\\src\\main\\scala\\CollisionDetector.scala 29:29]
  assign third_io_xPos = $signed(io_xPos) + $signed(_GEN_1204); // @[\\src\\main\\scala\\CollisionDetector.scala 30:28]
  assign third_io_yPos = $signed(io_yPos) + $signed(_GEN_1205); // @[\\src\\main\\scala\\CollisionDetector.scala 31:28]
  assign fourth_io_xPos = $signed(io_xPos) + $signed(_GEN_1206); // @[\\src\\main\\scala\\CollisionDetector.scala 32:29]
  assign fourth_io_yPos = $signed(io_yPos) + $signed(_GEN_1207); // @[\\src\\main\\scala\\CollisionDetector.scala 33:29]
endmodule
module PosToIndex(
  input  [10:0] io_xPos, // @[\\src\\main\\scala\\PosToIndex.scala 12:14]
  input  [9:0]  io_yPos, // @[\\src\\main\\scala\\PosToIndex.scala 12:14]
  output [10:0] io_index // @[\\src\\main\\scala\\PosToIndex.scala 12:14]
);
  wire [15:0] _io_index_T_1 = io_yPos * 6'h28; // @[\\src\\main\\scala\\PosToIndex.scala 18:30]
  wire [10:0] _io_index_T_2 = io_xPos; // @[\\src\\main\\scala\\PosToIndex.scala 18:47]
  wire [15:0] _GEN_0 = {{5'd0}, _io_index_T_2}; // @[\\src\\main\\scala\\PosToIndex.scala 18:37]
  wire [15:0] _io_index_T_4 = _io_index_T_1 + _GEN_0; // @[\\src\\main\\scala\\PosToIndex.scala 18:37]
  assign io_index = _io_index_T_4[10:0]; // @[\\src\\main\\scala\\PosToIndex.scala 18:12]
endmodule
module GameScreen(
  input        clock,
  input        reset,
  input        io_sw, // @[\\src\\main\\scala\\GameScreen.scala 7:14]
  output [9:0] io_viewBoxX, // @[\\src\\main\\scala\\GameScreen.scala 7:14]
  output [8:0] io_viewBoxY, // @[\\src\\main\\scala\\GameScreen.scala 7:14]
  output       io_staticScreen // @[\\src\\main\\scala\\GameScreen.scala 7:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] viewBoxXReg; // @[\\src\\main\\scala\\GameScreen.scala 17:28]
  reg [8:0] viewBoxYReg; // @[\\src\\main\\scala\\GameScreen.scala 18:28]
  reg [1:0] currentScreen; // @[\\src\\main\\scala\\GameScreen.scala 23:30]
  reg  static_; // @[\\src\\main\\scala\\GameScreen.scala 24:23]
  wire  _GEN_1 = 2'h2 == currentScreen | static_; // @[\\src\\main\\scala\\GameScreen.scala 28:24 43:14 24:23]
  wire  _GEN_6 = 2'h1 == currentScreen ? 1'h0 : _GEN_1; // @[\\src\\main\\scala\\GameScreen.scala 28:24 40:14]
  wire  _GEN_8 = 2'h0 == currentScreen | _GEN_6; // @[\\src\\main\\scala\\GameScreen.scala 28:24 33:14]
  assign io_viewBoxX = viewBoxXReg; // @[\\src\\main\\scala\\GameScreen.scala 19:15]
  assign io_viewBoxY = viewBoxYReg; // @[\\src\\main\\scala\\GameScreen.scala 20:15]
  assign io_staticScreen = static_; // @[\\src\\main\\scala\\GameScreen.scala 25:19]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GameScreen.scala 17:28]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GameScreen.scala 17:28]
    end else if (2'h0 == currentScreen) begin // @[\\src\\main\\scala\\GameScreen.scala 28:24]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GameScreen.scala 34:19]
    end else if (2'h1 == currentScreen) begin // @[\\src\\main\\scala\\GameScreen.scala 28:24]
      viewBoxXReg <= 10'h0; // @[\\src\\main\\scala\\GameScreen.scala 38:19]
    end else if (2'h2 == currentScreen) begin // @[\\src\\main\\scala\\GameScreen.scala 28:24]
      viewBoxXReg <= 10'h280; // @[\\src\\main\\scala\\GameScreen.scala 44:19]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameScreen.scala 18:28]
      viewBoxYReg <= 9'h0; // @[\\src\\main\\scala\\GameScreen.scala 18:28]
    end else if (2'h0 == currentScreen) begin // @[\\src\\main\\scala\\GameScreen.scala 28:24]
      viewBoxYReg <= 9'h1e0; // @[\\src\\main\\scala\\GameScreen.scala 35:19]
    end else if (2'h1 == currentScreen) begin // @[\\src\\main\\scala\\GameScreen.scala 28:24]
      viewBoxYReg <= 9'h0; // @[\\src\\main\\scala\\GameScreen.scala 39:19]
    end else if (2'h2 == currentScreen) begin // @[\\src\\main\\scala\\GameScreen.scala 28:24]
      viewBoxYReg <= 9'h1e0; // @[\\src\\main\\scala\\GameScreen.scala 45:19]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameScreen.scala 23:30]
      currentScreen <= 2'h0; // @[\\src\\main\\scala\\GameScreen.scala 23:30]
    end else if (2'h0 == currentScreen) begin // @[\\src\\main\\scala\\GameScreen.scala 28:24]
      if (io_sw) begin // @[\\src\\main\\scala\\GameScreen.scala 30:19]
        currentScreen <= 2'h1; // @[\\src\\main\\scala\\GameScreen.scala 31:23]
      end
    end
    static_ <= reset | _GEN_8; // @[\\src\\main\\scala\\GameScreen.scala 24:{23,23}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  viewBoxXReg = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  viewBoxYReg = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  currentScreen = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  static_ = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  input   io_increment, // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
  output  io_out_0, // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
  output  io_out_1, // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
  output  io_out_2 // @[src/main/scala/chisel3/util/random/PRNG.scala 42:22]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
  reg  state_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
  reg  state_2; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
  wire  _T = state_2 ^ state_1; // @[src/main/scala/chisel3/util/random/LFSR.scala 15:41]
  wire  _GEN_0 = io_increment ? _T : state_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 69:22 70:11 55:49]
  assign io_out_0 = state_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[src/main/scala/chisel3/util/random/PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _GEN_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:{49,49}]
    if (reset) begin // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
      state_1 <= 1'h0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
    end else if (io_increment) begin // @[src/main/scala/chisel3/util/random/PRNG.scala 69:22]
      state_1 <= state_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 70:11]
    end
    if (reset) begin // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
      state_2 <= 1'h0; // @[src/main/scala/chisel3/util/random/PRNG.scala 55:49]
    end else if (io_increment) begin // @[src/main/scala/chisel3/util/random/PRNG.scala 69:22]
      state_2 <= state_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 70:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BlockLogic(
  input  [1:0]  io_rotation, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  input  [10:0] io_xPos, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  input  [9:0]  io_yPos, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  input  [2:0]  io_sel, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_0, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_1, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_2, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_3, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_4, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_5, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_6, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_7, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_8, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_9, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_10, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_11, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_12, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_13, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_14, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_15, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_16, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_17, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_18, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_19, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_20, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_21, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_22, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_23, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_24, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_25, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_26, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [10:0] io_spriteXPosition_27, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_0, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_1, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_2, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_3, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_4, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_5, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_6, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_7, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_8, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_9, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_10, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_11, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_12, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_13, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_14, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_15, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_16, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_17, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_18, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_19, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_20, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_21, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_22, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_23, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_24, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_25, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_26, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [9:0]  io_spriteYPosition_27, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_0, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_1, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_2, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_3, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_4, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_5, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_6, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_7, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_8, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_9, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_10, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_11, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_12, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_13, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_14, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_15, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_16, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_17, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_18, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_19, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_20, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_21, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_22, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_23, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_24, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_25, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_26, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output        io_spriteVisible_27, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_activeOffsetX_0, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_activeOffsetX_1, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_activeOffsetX_2, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_activeOffsetX_3, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_activeOffsetY_0, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_activeOffsetY_1, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_activeOffsetY_2, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_activeOffsetY_3, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_nextOffsetX_0, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_nextOffsetX_1, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_nextOffsetX_2, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_nextOffsetX_3, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_nextOffsetY_0, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_nextOffsetY_1, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_nextOffsetY_2, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [3:0]  io_nextOffsetY_3, // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
  output [4:0]  io_tileNumber // @[\\src\\main\\scala\\BlockLogic.scala 5:14]
);
  wire [2:0] _T_1 = io_sel - 3'h1; // @[\\src\\main\\scala\\BlockLogic.scala 33:17]
  wire  _T_5 = io_rotation == 2'h0 | io_rotation == 2'h2; // @[\\src\\main\\scala\\BlockLogic.scala 36:32]
  wire [10:0] _io_spriteXPosition_0_T_2 = $signed(io_xPos) + 11'sh2; // @[\\src\\main\\scala\\BlockLogic.scala 39:45]
  wire [15:0] _io_spriteXPosition_0_T_3 = {$signed(_io_spriteXPosition_0_T_2), 5'h0}; // @[\\src\\main\\scala\\BlockLogic.scala 39:71]
  wire [9:0] _io_spriteYPosition_0_T_2 = $signed(io_yPos) + 10'sh1; // @[\\src\\main\\scala\\BlockLogic.scala 40:45]
  wire [14:0] _io_spriteYPosition_0_T_3 = {$signed(_io_spriteYPosition_0_T_2), 5'h0}; // @[\\src\\main\\scala\\BlockLogic.scala 40:71]
  wire [9:0] _io_spriteYPosition_1_T_2 = $signed(io_yPos) + 10'sh2; // @[\\src\\main\\scala\\BlockLogic.scala 40:45]
  wire [14:0] _io_spriteYPosition_1_T_3 = {$signed(_io_spriteYPosition_1_T_2), 5'h0}; // @[\\src\\main\\scala\\BlockLogic.scala 40:71]
  wire [10:0] _io_spriteXPosition_2_T_2 = $signed(io_xPos) + 11'sh3; // @[\\src\\main\\scala\\BlockLogic.scala 39:45]
  wire [15:0] _io_spriteXPosition_2_T_3 = {$signed(_io_spriteXPosition_2_T_2), 5'h0}; // @[\\src\\main\\scala\\BlockLogic.scala 39:71]
  wire [9:0] _io_spriteYPosition_3_T_2 = $signed(io_yPos) + 10'sh3; // @[\\src\\main\\scala\\BlockLogic.scala 40:45]
  wire [14:0] _io_spriteYPosition_3_T_3 = {$signed(_io_spriteYPosition_3_T_2), 5'h0}; // @[\\src\\main\\scala\\BlockLogic.scala 40:71]
  wire [10:0] _io_spriteXPosition_2_T_6 = $signed(io_xPos) + 11'sh1; // @[\\src\\main\\scala\\BlockLogic.scala 50:45]
  wire [15:0] _io_spriteXPosition_2_T_7 = {$signed(_io_spriteXPosition_2_T_6), 5'h0}; // @[\\src\\main\\scala\\BlockLogic.scala 50:72]
  wire [15:0] _GEN_1 = io_rotation == 2'h0 | io_rotation == 2'h2 ? $signed(_io_spriteXPosition_0_T_3) : $signed(
    _io_spriteXPosition_0_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 36:56 39:33 50:33]
  wire [14:0] _GEN_2 = io_rotation == 2'h0 | io_rotation == 2'h2 ? $signed(_io_spriteYPosition_0_T_3) : $signed(
    _io_spriteYPosition_0_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 36:56 40:33 51:33]
  wire [14:0] _GEN_4 = io_rotation == 2'h0 | io_rotation == 2'h2 ? $signed(_io_spriteYPosition_1_T_3) : $signed(
    _io_spriteYPosition_1_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 36:56 40:33 51:33]
  wire [15:0] _GEN_5 = io_rotation == 2'h0 | io_rotation == 2'h2 ? $signed(_io_spriteXPosition_2_T_3) : $signed(
    _io_spriteXPosition_2_T_7); // @[\\src\\main\\scala\\BlockLogic.scala 36:56 39:33 50:33]
  wire [15:0] _GEN_7 = io_rotation == 2'h0 | io_rotation == 2'h2 ? $signed(_io_spriteXPosition_2_T_3) : $signed(
    _io_spriteXPosition_2_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 36:56 39:33 50:33]
  wire [14:0] _GEN_8 = io_rotation == 2'h0 | io_rotation == 2'h2 ? $signed(_io_spriteYPosition_3_T_3) : $signed(
    _io_spriteYPosition_0_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 36:56 40:33 51:33]
  wire [3:0] _GEN_11 = io_rotation == 2'h0 | io_rotation == 2'h2 ? $signed(4'sh3) : $signed(4'sh1); // @[\\src\\main\\scala\\BlockLogic.scala 36:56 42:26 53:26]
  wire [3:0] _GEN_19 = io_rotation == 2'h0 | io_rotation == 2'h2 ? $signed(4'sh1) : $signed(4'sh3); // @[\\src\\main\\scala\\BlockLogic.scala 36:56 44:24 55:24]
  wire [15:0] _GEN_26 = _T_5 ? $signed(_io_spriteXPosition_2_T_3) : $signed(_io_spriteXPosition_0_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 63:56 66:33 77:33]
  wire [14:0] _GEN_27 = _T_5 ? $signed(_io_spriteYPosition_0_T_3) : $signed(_io_spriteYPosition_3_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 63:56 67:33 78:33]
  wire [15:0] _GEN_30 = _T_5 ? $signed(_io_spriteXPosition_0_T_3) : $signed(_io_spriteXPosition_2_T_7); // @[\\src\\main\\scala\\BlockLogic.scala 63:56 66:33 77:33]
  wire [15:0] _GEN_32 = _T_5 ? $signed(_io_spriteXPosition_0_T_3) : $signed(_io_spriteXPosition_2_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 63:56 66:33 77:33]
  wire [14:0] _GEN_33 = _T_5 ? $signed(_io_spriteYPosition_3_T_3) : $signed(_io_spriteYPosition_3_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 63:56 67:33 78:33]
  wire [3:0] _GEN_34 = _T_5 ? $signed(4'sh3) : $signed(4'sh2); // @[\\src\\main\\scala\\BlockLogic.scala 63:56 69:26 80:26]
  wire [3:0] _GEN_36 = _T_5 ? $signed(4'sh2) : $signed(4'sh1); // @[\\src\\main\\scala\\BlockLogic.scala 63:56 69:26 80:26]
  wire [3:0] _GEN_37 = _T_5 ? $signed(4'sh2) : $signed(4'sh3); // @[\\src\\main\\scala\\BlockLogic.scala 63:56 69:26 80:26]
  wire [3:0] _GEN_44 = _T_5 ? $signed(4'sh1) : $signed(4'sh2); // @[\\src\\main\\scala\\BlockLogic.scala 63:56 71:24 82:24]
  wire [11:0] _io_spriteXPosition_12_T = {{1{io_xPos[10]}},io_xPos}; // @[\\src\\main\\scala\\BlockLogic.scala 106:45]
  wire [10:0] _io_spriteXPosition_12_T_2 = _io_spriteXPosition_12_T[10:0]; // @[\\src\\main\\scala\\BlockLogic.scala 106:45]
  wire [15:0] _io_spriteXPosition_12_T_3 = {$signed(_io_spriteXPosition_12_T_2), 5'h0}; // @[\\src\\main\\scala\\BlockLogic.scala 106:77]
  wire [10:0] _io_spriteYPosition_12_T_4 = {{1{io_yPos[9]}},io_yPos}; // @[\\src\\main\\scala\\BlockLogic.scala 117:45]
  wire [9:0] _io_spriteYPosition_12_T_6 = _io_spriteYPosition_12_T_4[9:0]; // @[\\src\\main\\scala\\BlockLogic.scala 117:45]
  wire [14:0] _io_spriteYPosition_12_T_7 = {$signed(_io_spriteYPosition_12_T_6), 5'h0}; // @[\\src\\main\\scala\\BlockLogic.scala 117:78]
  wire [15:0] _GEN_51 = _T_5 ? $signed(_io_spriteXPosition_12_T_3) : $signed(_io_spriteXPosition_0_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 103:56 106:33 116:33]
  wire [14:0] _GEN_52 = _T_5 ? $signed(_io_spriteYPosition_1_T_3) : $signed(_io_spriteYPosition_12_T_7); // @[\\src\\main\\scala\\BlockLogic.scala 103:56 107:33 117:33]
  wire [15:0] _GEN_53 = _T_5 ? $signed(_io_spriteXPosition_2_T_7) : $signed(_io_spriteXPosition_0_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 103:56 106:33 116:33]
  wire [14:0] _GEN_54 = _T_5 ? $signed(_io_spriteYPosition_1_T_3) : $signed(_io_spriteYPosition_0_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 103:56 107:33 117:33]
  wire [14:0] _GEN_58 = _T_5 ? $signed(_io_spriteYPosition_1_T_3) : $signed(_io_spriteYPosition_3_T_3); // @[\\src\\main\\scala\\BlockLogic.scala 103:56 107:33 117:33]
  wire [3:0] _GEN_59 = _T_5 ? $signed(4'sh0) : $signed(4'sh2); // @[\\src\\main\\scala\\BlockLogic.scala 103:56 109:26 119:26]
  wire [3:0] _GEN_63 = _T_5 ? $signed(4'sh2) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 103:56 110:26 120:26]
  wire  _T_16 = 2'h0 == io_rotation; // @[\\src\\main\\scala\\BlockLogic.scala 129:26]
  wire  _T_17 = 2'h1 == io_rotation; // @[\\src\\main\\scala\\BlockLogic.scala 129:26]
  wire  _T_18 = 2'h2 == io_rotation; // @[\\src\\main\\scala\\BlockLogic.scala 129:26]
  wire  _T_19 = 2'h3 == io_rotation; // @[\\src\\main\\scala\\BlockLogic.scala 129:26]
  wire [15:0] _GEN_76 = 2'h3 == io_rotation ? $signed(_io_spriteXPosition_2_T_3) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 169:35 20:22]
  wire [14:0] _GEN_77 = 2'h3 == io_rotation ? $signed(_io_spriteYPosition_3_T_3) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 170:35 21:22]
  wire [14:0] _GEN_79 = 2'h3 == io_rotation ? $signed(_io_spriteYPosition_1_T_3) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 170:35 21:22]
  wire [14:0] _GEN_81 = 2'h3 == io_rotation ? $signed(_io_spriteYPosition_0_T_3) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 170:35 21:22]
  wire [15:0] _GEN_82 = 2'h3 == io_rotation ? $signed(_io_spriteXPosition_0_T_3) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 169:35 20:22]
  wire [3:0] _GEN_84 = 2'h3 == io_rotation ? $signed(4'sh3) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 172:28 23:20]
  wire [3:0] _GEN_87 = 2'h3 == io_rotation ? $signed(4'sh2) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 172:28 23:20]
  wire [3:0] _GEN_90 = 2'h3 == io_rotation ? $signed(4'sh1) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 173:28 24:20]
  wire  _GEN_100 = 2'h2 == io_rotation | 2'h3 == io_rotation; // @[\\src\\main\\scala\\BlockLogic.scala 129:26 156:33]
  wire [15:0] _GEN_101 = 2'h2 == io_rotation ? $signed(_io_spriteXPosition_2_T_7) : $signed(_GEN_76); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 157:35]
  wire [14:0] _GEN_102 = 2'h2 == io_rotation ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_77); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 158:35]
  wire [15:0] _GEN_103 = 2'h2 == io_rotation ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_76); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 157:35]
  wire [14:0] _GEN_104 = 2'h2 == io_rotation ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_79); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 158:35]
  wire [15:0] _GEN_105 = 2'h2 == io_rotation ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_76); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 157:35]
  wire [14:0] _GEN_106 = 2'h2 == io_rotation ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_81); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 158:35]
  wire [15:0] _GEN_107 = 2'h2 == io_rotation ? $signed(_io_spriteXPosition_2_T_7) : $signed(_GEN_82); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 157:35]
  wire [14:0] _GEN_108 = 2'h2 == io_rotation ? $signed(_io_spriteYPosition_3_T_3) : $signed(_GEN_81); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 158:35]
  wire [3:0] _GEN_109 = 2'h2 == io_rotation ? $signed(4'sh1) : $signed(_GEN_84); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 160:28]
  wire [3:0] _GEN_110 = 2'h2 == io_rotation ? $signed(4'sh2) : $signed(_GEN_84); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 160:28]
  wire [3:0] _GEN_111 = 2'h2 == io_rotation ? $signed(4'sh3) : $signed(_GEN_84); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 160:28]
  wire [3:0] _GEN_112 = 2'h2 == io_rotation ? $signed(4'sh1) : $signed(_GEN_87); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 160:28]
  wire [3:0] _GEN_114 = 2'h2 == io_rotation ? $signed(4'sh2) : $signed(_GEN_87); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 161:28]
  wire [3:0] _GEN_115 = 2'h2 == io_rotation ? $signed(4'sh2) : $signed(_GEN_90); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 161:28]
  wire [3:0] _GEN_116 = 2'h2 == io_rotation ? $signed(4'sh3) : $signed(_GEN_90); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 161:28]
  wire [3:0] _GEN_118 = 2'h2 == io_rotation ? $signed(4'sh3) : $signed(_GEN_87); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 162:26]
  wire [3:0] _GEN_124 = 2'h2 == io_rotation ? $signed(4'sh1) : $signed(_GEN_90); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 163:26]
  wire  _GEN_125 = 2'h1 == io_rotation | _GEN_100; // @[\\src\\main\\scala\\BlockLogic.scala 129:26 144:33]
  wire [15:0] _GEN_126 = 2'h1 == io_rotation ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_101); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 145:35]
  wire [14:0] _GEN_127 = 2'h1 == io_rotation ? $signed(_io_spriteYPosition_0_T_3) : $signed(_GEN_102); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 146:35]
  wire [15:0] _GEN_128 = 2'h1 == io_rotation ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_103); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 145:35]
  wire [14:0] _GEN_129 = 2'h1 == io_rotation ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_104); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 146:35]
  wire [15:0] _GEN_130 = 2'h1 == io_rotation ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_105); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 145:35]
  wire [14:0] _GEN_131 = 2'h1 == io_rotation ? $signed(_io_spriteYPosition_3_T_3) : $signed(_GEN_106); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 146:35]
  wire [15:0] _GEN_132 = 2'h1 == io_rotation ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_107); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 145:35]
  wire [14:0] _GEN_133 = 2'h1 == io_rotation ? $signed(_io_spriteYPosition_3_T_3) : $signed(_GEN_108); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 146:35]
  wire [3:0] _GEN_134 = 2'h1 == io_rotation ? $signed(4'sh2) : $signed(_GEN_109); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 148:28]
  wire [3:0] _GEN_135 = 2'h1 == io_rotation ? $signed(4'sh2) : $signed(_GEN_110); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 148:28]
  wire [3:0] _GEN_136 = 2'h1 == io_rotation ? $signed(4'sh2) : $signed(_GEN_111); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 148:28]
  wire [3:0] _GEN_137 = 2'h1 == io_rotation ? $signed(4'sh3) : $signed(_GEN_112); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 148:28]
  wire [3:0] _GEN_138 = 2'h1 == io_rotation ? $signed(4'sh1) : $signed(_GEN_110); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 149:28]
  wire [3:0] _GEN_139 = 2'h1 == io_rotation ? $signed(4'sh2) : $signed(_GEN_114); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 149:28]
  wire [3:0] _GEN_140 = 2'h1 == io_rotation ? $signed(4'sh3) : $signed(_GEN_115); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 149:28]
  wire [3:0] _GEN_141 = 2'h1 == io_rotation ? $signed(4'sh3) : $signed(_GEN_116); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 149:28]
  wire [3:0] _GEN_142 = 2'h1 == io_rotation ? $signed(4'sh1) : $signed(_GEN_116); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 150:26]
  wire [3:0] _GEN_143 = 2'h1 == io_rotation ? $signed(4'sh2) : $signed(_GEN_118); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 150:26]
  wire [3:0] _GEN_144 = 2'h1 == io_rotation ? $signed(4'sh3) : $signed(_GEN_111); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 150:26]
  wire [3:0] _GEN_148 = 2'h1 == io_rotation ? $signed(4'sh2) : $signed(_GEN_112); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 151:26]
  wire [3:0] _GEN_149 = 2'h1 == io_rotation ? $signed(4'sh3) : $signed(_GEN_124); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 151:26]
  wire  _GEN_150 = 2'h0 == io_rotation | _GEN_125; // @[\\src\\main\\scala\\BlockLogic.scala 129:26 132:33]
  wire [15:0] _GEN_151 = 2'h0 == io_rotation ? $signed(_io_spriteXPosition_2_T_7) : $signed(_GEN_126); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 133:35]
  wire [14:0] _GEN_152 = 2'h0 == io_rotation ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_127); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 134:35]
  wire [15:0] _GEN_153 = 2'h0 == io_rotation ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_128); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 133:35]
  wire [14:0] _GEN_154 = 2'h0 == io_rotation ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_129); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 134:35]
  wire [15:0] _GEN_155 = 2'h0 == io_rotation ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_130); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 133:35]
  wire [14:0] _GEN_156 = 2'h0 == io_rotation ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_131); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 134:35]
  wire [15:0] _GEN_157 = 2'h0 == io_rotation ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_132); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 133:35]
  wire [14:0] _GEN_158 = 2'h0 == io_rotation ? $signed(_io_spriteYPosition_0_T_3) : $signed(_GEN_133); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 134:35]
  wire [3:0] _GEN_159 = 2'h0 == io_rotation ? $signed(4'sh1) : $signed(_GEN_134); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 136:28]
  wire [3:0] _GEN_160 = 2'h0 == io_rotation ? $signed(4'sh2) : $signed(_GEN_135); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 136:28]
  wire [3:0] _GEN_161 = 2'h0 == io_rotation ? $signed(4'sh3) : $signed(_GEN_136); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 136:28]
  wire [3:0] _GEN_162 = 2'h0 == io_rotation ? $signed(4'sh3) : $signed(_GEN_137); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 136:28]
  wire [3:0] _GEN_163 = 2'h0 == io_rotation ? $signed(4'sh2) : $signed(_GEN_138); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 137:28]
  wire [3:0] _GEN_164 = 2'h0 == io_rotation ? $signed(4'sh2) : $signed(_GEN_139); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 137:28]
  wire [3:0] _GEN_165 = 2'h0 == io_rotation ? $signed(4'sh2) : $signed(_GEN_140); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 137:28]
  wire [3:0] _GEN_166 = 2'h0 == io_rotation ? $signed(4'sh1) : $signed(_GEN_141); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 137:28]
  wire [3:0] _GEN_167 = 2'h0 == io_rotation ? $signed(4'sh2) : $signed(_GEN_142); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 138:26]
  wire [3:0] _GEN_168 = 2'h0 == io_rotation ? $signed(4'sh2) : $signed(_GEN_143); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 138:26]
  wire [3:0] _GEN_169 = 2'h0 == io_rotation ? $signed(4'sh2) : $signed(_GEN_144); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 138:26]
  wire [3:0] _GEN_170 = 2'h0 == io_rotation ? $signed(4'sh3) : $signed(_GEN_138); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 138:26]
  wire [3:0] _GEN_171 = 2'h0 == io_rotation ? $signed(4'sh1) : $signed(_GEN_143); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 139:26]
  wire [3:0] _GEN_173 = 2'h0 == io_rotation ? $signed(4'sh3) : $signed(_GEN_148); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 139:26]
  wire [3:0] _GEN_174 = 2'h0 == io_rotation ? $signed(4'sh3) : $signed(_GEN_149); // @[\\src\\main\\scala\\BlockLogic.scala 129:26 139:26]
  wire [15:0] _GEN_203 = _T_18 ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_82); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 210:35]
  wire [15:0] _GEN_205 = _T_18 ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_82); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 210:35]
  wire [14:0] _GEN_208 = _T_18 ? $signed(_io_spriteYPosition_0_T_3) : $signed(_GEN_77); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 211:35]
  wire [15:0] _GEN_228 = _T_17 ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_203); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 198:35]
  wire [15:0] _GEN_230 = _T_17 ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_205); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 198:35]
  wire [14:0] _GEN_233 = _T_17 ? $signed(_io_spriteYPosition_0_T_3) : $signed(_GEN_208); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 199:35]
  wire [3:0] _GEN_235 = _T_17 ? $signed(4'sh3) : $signed(_GEN_114); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 201:28]
  wire [3:0] _GEN_236 = _T_17 ? $signed(4'sh3) : $signed(_GEN_118); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 201:28]
  wire [3:0] _GEN_241 = _T_17 ? $signed(4'sh1) : $signed(_GEN_109); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 202:28]
  wire [3:0] _GEN_244 = _T_17 ? $signed(4'sh3) : $signed(_GEN_110); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 203:26]
  wire [3:0] _GEN_249 = _T_17 ? $signed(4'sh1) : $signed(_GEN_111); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 204:26]
  wire [15:0] _GEN_253 = _T_16 ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_228); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 186:35]
  wire [15:0] _GEN_255 = _T_16 ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_230); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 186:35]
  wire [14:0] _GEN_258 = _T_16 ? $signed(_io_spriteYPosition_3_T_3) : $signed(_GEN_233); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 187:35]
  wire [3:0] _GEN_260 = _T_16 ? $signed(4'sh2) : $signed(_GEN_235); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 189:28]
  wire [3:0] _GEN_261 = _T_16 ? $signed(4'sh3) : $signed(_GEN_236); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 189:28]
  wire [3:0] _GEN_266 = _T_16 ? $signed(4'sh3) : $signed(_GEN_241); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 190:28]
  wire [3:0] _GEN_268 = _T_16 ? $signed(4'sh3) : $signed(_GEN_139); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 191:26]
  wire [3:0] _GEN_269 = _T_16 ? $signed(4'sh3) : $signed(_GEN_244); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 191:26]
  wire [3:0] _GEN_274 = _T_16 ? $signed(4'sh1) : $signed(_GEN_249); // @[\\src\\main\\scala\\BlockLogic.scala 182:26 192:26]
  wire [15:0] _GEN_280 = _T_19 ? $signed(_io_spriteXPosition_2_T_7) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 234:27 273:35]
  wire [14:0] _GEN_302 = _T_18 ? $signed(_io_spriteYPosition_3_T_3) : $signed(_GEN_77); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 263:35]
  wire [15:0] _GEN_305 = _T_18 ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_280); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 262:35]
  wire [14:0] _GEN_308 = _T_18 ? $signed(_io_spriteYPosition_0_T_3) : $signed(_GEN_79); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 263:35]
  wire [15:0] _GEN_326 = _T_17 ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_203); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 250:35]
  wire [14:0] _GEN_327 = _T_17 ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_302); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 251:35]
  wire [15:0] _GEN_328 = _T_17 ? $signed(_io_spriteXPosition_2_T_7) : $signed(_GEN_203); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 250:35]
  wire [15:0] _GEN_330 = _T_17 ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_305); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 250:35]
  wire [14:0] _GEN_331 = _T_17 ? $signed(_io_spriteYPosition_0_T_3) : $signed(_GEN_104); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 251:35]
  wire [15:0] _GEN_332 = _T_17 ? $signed(_io_spriteXPosition_2_T_3) : $signed(_GEN_103); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 250:35]
  wire [14:0] _GEN_333 = _T_17 ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_308); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 251:35]
  wire [3:0] _GEN_335 = _T_17 ? $signed(4'sh1) : $signed(_GEN_114); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 253:28]
  wire [3:0] _GEN_336 = _T_17 ? $signed(4'sh2) : $signed(_GEN_116); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 253:28]
  wire [3:0] _GEN_349 = _T_17 ? $signed(4'sh1) : $signed(_GEN_115); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 256:26]
  wire [15:0] _GEN_351 = _T_16 ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_326); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 238:35]
  wire [14:0] _GEN_352 = _T_16 ? $signed(_io_spriteYPosition_3_T_3) : $signed(_GEN_327); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 239:35]
  wire [15:0] _GEN_353 = _T_16 ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_328); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 238:35]
  wire [15:0] _GEN_355 = _T_16 ? $signed(_io_spriteXPosition_2_T_7) : $signed(_GEN_330); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 238:35]
  wire [14:0] _GEN_356 = _T_16 ? $signed(_io_spriteYPosition_1_T_3) : $signed(_GEN_331); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 239:35]
  wire [15:0] _GEN_357 = _T_16 ? $signed(_io_spriteXPosition_0_T_3) : $signed(_GEN_332); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 238:35]
  wire [14:0] _GEN_358 = _T_16 ? $signed(_io_spriteYPosition_0_T_3) : $signed(_GEN_333); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 239:35]
  wire [3:0] _GEN_360 = _T_16 ? $signed(4'sh2) : $signed(_GEN_335); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 241:28]
  wire [3:0] _GEN_361 = _T_16 ? $signed(4'sh1) : $signed(_GEN_336); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 241:28]
  wire [3:0] _GEN_362 = _T_16 ? $signed(4'sh2) : $signed(_GEN_244); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 241:28]
  wire [3:0] _GEN_366 = _T_16 ? $signed(4'sh1) : $signed(_GEN_148); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 242:28]
  wire [3:0] _GEN_368 = _T_16 ? $signed(4'sh1) : $signed(_GEN_139); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 243:26]
  wire [3:0] _GEN_369 = _T_16 ? $signed(4'sh2) : $signed(_GEN_149); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 243:26]
  wire [3:0] _GEN_370 = _T_16 ? $signed(4'sh3) : $signed(_GEN_143); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 243:26]
  wire [3:0] _GEN_374 = _T_16 ? $signed(4'sh2) : $signed(_GEN_349); // @[\\src\\main\\scala\\BlockLogic.scala 234:27 244:26]
  wire [15:0] _GEN_376 = 3'h6 == _T_1 ? $signed(_GEN_351) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_377 = 3'h6 == _T_1 ? $signed(_GEN_352) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_378 = 3'h6 == _T_1 ? $signed(_GEN_353) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_379 = 3'h6 == _T_1 ? $signed(_GEN_154) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_380 = 3'h6 == _T_1 ? $signed(_GEN_355) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_381 = 3'h6 == _T_1 ? $signed(_GEN_356) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_382 = 3'h6 == _T_1 ? $signed(_GEN_357) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_383 = 3'h6 == _T_1 ? $signed(_GEN_358) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [3:0] _GEN_384 = 3'h6 == _T_1 ? $signed(_GEN_164) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 23:20 33:23]
  wire [3:0] _GEN_385 = 3'h6 == _T_1 ? $signed(_GEN_360) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 23:20 33:23]
  wire [3:0] _GEN_386 = 3'h6 == _T_1 ? $signed(_GEN_361) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 23:20 33:23]
  wire [3:0] _GEN_387 = 3'h6 == _T_1 ? $signed(_GEN_362) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 23:20 33:23]
  wire [3:0] _GEN_388 = 3'h6 == _T_1 ? $signed(_GEN_161) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 24:20 33:23]
  wire [3:0] _GEN_391 = 3'h6 == _T_1 ? $signed(_GEN_366) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 24:20 33:23]
  wire [3:0] _GEN_393 = 3'h6 == _T_1 ? $signed(_GEN_368) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 25:18 33:23]
  wire [3:0] _GEN_394 = 3'h6 == _T_1 ? $signed(_GEN_369) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 25:18 33:23]
  wire [3:0] _GEN_395 = 3'h6 == _T_1 ? $signed(_GEN_370) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 25:18 33:23]
  wire [3:0] _GEN_396 = 3'h6 == _T_1 ? $signed(_GEN_169) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 26:18 33:23]
  wire [3:0] _GEN_399 = 3'h6 == _T_1 ? $signed(_GEN_374) : $signed(4'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 26:18 33:23]
  wire [4:0] _GEN_400 = 3'h6 == _T_1 ? 5'h1b : 5'h0; // @[\\src\\main\\scala\\BlockLogic.scala 27:17 282:21 33:23]
  wire [15:0] _GEN_402 = 3'h5 == _T_1 ? $signed(_GEN_151) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_403 = 3'h5 == _T_1 ? $signed(_GEN_156) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_404 = 3'h5 == _T_1 ? $signed(_GEN_253) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_406 = 3'h5 == _T_1 ? $signed(_GEN_255) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_407 = 3'h5 == _T_1 ? $signed(_GEN_154) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_408 = 3'h5 == _T_1 ? $signed(_GEN_157) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_409 = 3'h5 == _T_1 ? $signed(_GEN_258) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [3:0] _GEN_410 = 3'h5 == _T_1 ? $signed(_GEN_159) : $signed(_GEN_384); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_411 = 3'h5 == _T_1 ? $signed(_GEN_260) : $signed(_GEN_385); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_412 = 3'h5 == _T_1 ? $signed(_GEN_261) : $signed(_GEN_386); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_413 = 3'h5 == _T_1 ? $signed(_GEN_162) : $signed(_GEN_387); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_414 = 3'h5 == _T_1 ? $signed(_GEN_165) : $signed(_GEN_388); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_415 = 3'h5 == _T_1 ? $signed(_GEN_165) : $signed(_GEN_384); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_416 = 3'h5 == _T_1 ? $signed(_GEN_164) : $signed(_GEN_385); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_417 = 3'h5 == _T_1 ? $signed(_GEN_266) : $signed(_GEN_391); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_418 = 3'h5 == _T_1 ? $signed(_GEN_167) : $signed(_GEN_384); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_419 = 3'h5 == _T_1 ? $signed(_GEN_268) : $signed(_GEN_393); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_420 = 3'h5 == _T_1 ? $signed(_GEN_269) : $signed(_GEN_394); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_421 = 3'h5 == _T_1 ? $signed(_GEN_170) : $signed(_GEN_395); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_422 = 3'h5 == _T_1 ? $signed(_GEN_173) : $signed(_GEN_396); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_423 = 3'h5 == _T_1 ? $signed(_GEN_173) : $signed(_GEN_384); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_424 = 3'h5 == _T_1 ? $signed(_GEN_164) : $signed(_GEN_393); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_425 = 3'h5 == _T_1 ? $signed(_GEN_274) : $signed(_GEN_399); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [4:0] _GEN_426 = 3'h5 == _T_1 ? 5'h1a : _GEN_400; // @[\\src\\main\\scala\\BlockLogic.scala 231:21 33:23]
  wire  _GEN_427 = 3'h5 == _T_1 ? 1'h0 : 3'h6 == _T_1 & _GEN_150; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_428 = 3'h5 == _T_1 ? $signed(16'sh0) : $signed(_GEN_376); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_429 = 3'h5 == _T_1 ? $signed(15'sh0) : $signed(_GEN_377); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_430 = 3'h5 == _T_1 ? $signed(16'sh0) : $signed(_GEN_378); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_431 = 3'h5 == _T_1 ? $signed(15'sh0) : $signed(_GEN_379); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_432 = 3'h5 == _T_1 ? $signed(16'sh0) : $signed(_GEN_380); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_433 = 3'h5 == _T_1 ? $signed(15'sh0) : $signed(_GEN_381); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_434 = 3'h5 == _T_1 ? $signed(16'sh0) : $signed(_GEN_382); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_435 = 3'h5 == _T_1 ? $signed(15'sh0) : $signed(_GEN_383); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_437 = 3'h4 == _T_1 ? $signed(_GEN_151) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_438 = 3'h4 == _T_1 ? $signed(_GEN_152) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_439 = 3'h4 == _T_1 ? $signed(_GEN_153) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_440 = 3'h4 == _T_1 ? $signed(_GEN_154) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_441 = 3'h4 == _T_1 ? $signed(_GEN_155) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_442 = 3'h4 == _T_1 ? $signed(_GEN_156) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_443 = 3'h4 == _T_1 ? $signed(_GEN_157) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_444 = 3'h4 == _T_1 ? $signed(_GEN_158) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [3:0] _GEN_445 = 3'h4 == _T_1 ? $signed(_GEN_159) : $signed(_GEN_410); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_446 = 3'h4 == _T_1 ? $signed(_GEN_160) : $signed(_GEN_411); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_447 = 3'h4 == _T_1 ? $signed(_GEN_161) : $signed(_GEN_412); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_448 = 3'h4 == _T_1 ? $signed(_GEN_162) : $signed(_GEN_413); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_449 = 3'h4 == _T_1 ? $signed(_GEN_163) : $signed(_GEN_414); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_450 = 3'h4 == _T_1 ? $signed(_GEN_164) : $signed(_GEN_415); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_451 = 3'h4 == _T_1 ? $signed(_GEN_165) : $signed(_GEN_416); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_452 = 3'h4 == _T_1 ? $signed(_GEN_166) : $signed(_GEN_417); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_453 = 3'h4 == _T_1 ? $signed(_GEN_167) : $signed(_GEN_418); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_454 = 3'h4 == _T_1 ? $signed(_GEN_168) : $signed(_GEN_419); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_455 = 3'h4 == _T_1 ? $signed(_GEN_169) : $signed(_GEN_420); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_456 = 3'h4 == _T_1 ? $signed(_GEN_170) : $signed(_GEN_421); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_457 = 3'h4 == _T_1 ? $signed(_GEN_171) : $signed(_GEN_422); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_458 = 3'h4 == _T_1 ? $signed(_GEN_164) : $signed(_GEN_423); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_459 = 3'h4 == _T_1 ? $signed(_GEN_173) : $signed(_GEN_424); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_460 = 3'h4 == _T_1 ? $signed(_GEN_174) : $signed(_GEN_425); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [4:0] _GEN_461 = 3'h4 == _T_1 ? 5'h19 : _GEN_426; // @[\\src\\main\\scala\\BlockLogic.scala 179:21 33:23]
  wire  _GEN_462 = 3'h4 == _T_1 ? 1'h0 : 3'h5 == _T_1 & _GEN_150; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_463 = 3'h4 == _T_1 ? $signed(16'sh0) : $signed(_GEN_402); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_464 = 3'h4 == _T_1 ? $signed(15'sh0) : $signed(_GEN_403); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_465 = 3'h4 == _T_1 ? $signed(16'sh0) : $signed(_GEN_404); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_467 = 3'h4 == _T_1 ? $signed(16'sh0) : $signed(_GEN_406); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_468 = 3'h4 == _T_1 ? $signed(15'sh0) : $signed(_GEN_407); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_469 = 3'h4 == _T_1 ? $signed(16'sh0) : $signed(_GEN_408); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_470 = 3'h4 == _T_1 ? $signed(15'sh0) : $signed(_GEN_409); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire  _GEN_471 = 3'h4 == _T_1 ? 1'h0 : _GEN_427; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_472 = 3'h4 == _T_1 ? $signed(16'sh0) : $signed(_GEN_428); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_473 = 3'h4 == _T_1 ? $signed(15'sh0) : $signed(_GEN_429); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_474 = 3'h4 == _T_1 ? $signed(16'sh0) : $signed(_GEN_430); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_475 = 3'h4 == _T_1 ? $signed(15'sh0) : $signed(_GEN_431); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_476 = 3'h4 == _T_1 ? $signed(16'sh0) : $signed(_GEN_432); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_477 = 3'h4 == _T_1 ? $signed(15'sh0) : $signed(_GEN_433); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_478 = 3'h4 == _T_1 ? $signed(16'sh0) : $signed(_GEN_434); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_479 = 3'h4 == _T_1 ? $signed(15'sh0) : $signed(_GEN_435); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_481 = 3'h3 == _T_1 ? $signed(_GEN_51) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_482 = 3'h3 == _T_1 ? $signed(_GEN_52) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_483 = 3'h3 == _T_1 ? $signed(_GEN_53) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_484 = 3'h3 == _T_1 ? $signed(_GEN_54) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_485 = 3'h3 == _T_1 ? $signed(_GEN_1) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_486 = 3'h3 == _T_1 ? $signed(_GEN_4) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_487 = 3'h3 == _T_1 ? $signed(_GEN_26) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_488 = 3'h3 == _T_1 ? $signed(_GEN_58) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [3:0] _GEN_489 = 3'h3 == _T_1 ? $signed(_GEN_59) : $signed(_GEN_445); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_490 = 3'h3 == _T_1 ? $signed(_GEN_44) : $signed(_GEN_446); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_491 = 3'h3 == _T_1 ? $signed(4'sh2) : $signed(_GEN_447); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_492 = 3'h3 == _T_1 ? $signed(_GEN_34) : $signed(_GEN_448); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_493 = 3'h3 == _T_1 ? $signed(_GEN_63) : $signed(_GEN_449); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_494 = 3'h3 == _T_1 ? $signed(_GEN_36) : $signed(_GEN_450); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_495 = 3'h3 == _T_1 ? $signed(4'sh2) : $signed(_GEN_451); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_496 = 3'h3 == _T_1 ? $signed(_GEN_37) : $signed(_GEN_452); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_497 = 3'h3 == _T_1 ? $signed(_GEN_63) : $signed(_GEN_453); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_498 = 3'h3 == _T_1 ? $signed(_GEN_36) : $signed(_GEN_454); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_499 = 3'h3 == _T_1 ? $signed(4'sh2) : $signed(_GEN_455); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_500 = 3'h3 == _T_1 ? $signed(_GEN_37) : $signed(_GEN_456); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_501 = 3'h3 == _T_1 ? $signed(_GEN_59) : $signed(_GEN_457); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_502 = 3'h3 == _T_1 ? $signed(_GEN_44) : $signed(_GEN_458); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_503 = 3'h3 == _T_1 ? $signed(4'sh2) : $signed(_GEN_459); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_504 = 3'h3 == _T_1 ? $signed(_GEN_34) : $signed(_GEN_460); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [4:0] _GEN_505 = 3'h3 == _T_1 ? 5'h18 : _GEN_461; // @[\\src\\main\\scala\\BlockLogic.scala 125:21 33:23]
  wire  _GEN_506 = 3'h3 == _T_1 ? 1'h0 : 3'h4 == _T_1 & _GEN_150; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_507 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_437); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_508 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_438); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_509 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_439); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_510 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_440); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_511 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_441); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_512 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_442); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_513 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_443); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_514 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_444); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire  _GEN_515 = 3'h3 == _T_1 ? 1'h0 : _GEN_462; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_516 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_463); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_517 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_464); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_518 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_465); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_520 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_467); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_521 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_468); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_522 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_469); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_523 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_470); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire  _GEN_524 = 3'h3 == _T_1 ? 1'h0 : _GEN_471; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_525 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_472); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_526 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_473); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_527 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_474); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_528 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_475); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_529 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_476); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_530 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_477); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_531 = 3'h3 == _T_1 ? $signed(16'sh0) : $signed(_GEN_478); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_532 = 3'h3 == _T_1 ? $signed(15'sh0) : $signed(_GEN_479); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_534 = 3'h2 == _T_1 ? $signed(_io_spriteXPosition_0_T_3) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23 92:31]
  wire [14:0] _GEN_535 = 3'h2 == _T_1 ? $signed(_io_spriteYPosition_0_T_3) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23 93:31]
  wire [14:0] _GEN_537 = 3'h2 == _T_1 ? $signed(_io_spriteYPosition_1_T_3) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23 93:31]
  wire [15:0] _GEN_538 = 3'h2 == _T_1 ? $signed(_io_spriteXPosition_2_T_3) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23 92:31]
  wire [3:0] _GEN_542 = 3'h2 == _T_1 ? $signed(4'sh2) : $signed(_GEN_489); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 95:24]
  wire [3:0] _GEN_543 = 3'h2 == _T_1 ? $signed(4'sh2) : $signed(_GEN_490); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 95:24]
  wire [3:0] _GEN_544 = 3'h2 == _T_1 ? $signed(4'sh3) : $signed(_GEN_491); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 95:24]
  wire [3:0] _GEN_545 = 3'h2 == _T_1 ? $signed(4'sh3) : $signed(_GEN_492); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 95:24]
  wire [3:0] _GEN_546 = 3'h2 == _T_1 ? $signed(4'sh1) : $signed(_GEN_493); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 96:24]
  wire [3:0] _GEN_547 = 3'h2 == _T_1 ? $signed(4'sh2) : $signed(_GEN_494); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 96:24]
  wire [3:0] _GEN_548 = 3'h2 == _T_1 ? $signed(4'sh1) : $signed(_GEN_495); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 96:24]
  wire [3:0] _GEN_549 = 3'h2 == _T_1 ? $signed(4'sh2) : $signed(_GEN_496); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 96:24]
  wire [3:0] _GEN_550 = 3'h2 == _T_1 ? $signed(4'sh2) : $signed(_GEN_497); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 97:22]
  wire [3:0] _GEN_551 = 3'h2 == _T_1 ? $signed(4'sh2) : $signed(_GEN_498); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 97:22]
  wire [3:0] _GEN_552 = 3'h2 == _T_1 ? $signed(4'sh3) : $signed(_GEN_499); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 97:22]
  wire [3:0] _GEN_553 = 3'h2 == _T_1 ? $signed(4'sh3) : $signed(_GEN_500); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 97:22]
  wire [3:0] _GEN_554 = 3'h2 == _T_1 ? $signed(4'sh1) : $signed(_GEN_501); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 98:22]
  wire [3:0] _GEN_555 = 3'h2 == _T_1 ? $signed(4'sh2) : $signed(_GEN_502); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 98:22]
  wire [3:0] _GEN_556 = 3'h2 == _T_1 ? $signed(4'sh1) : $signed(_GEN_503); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 98:22]
  wire [3:0] _GEN_557 = 3'h2 == _T_1 ? $signed(4'sh2) : $signed(_GEN_504); // @[\\src\\main\\scala\\BlockLogic.scala 33:23 98:22]
  wire [4:0] _GEN_558 = 3'h2 == _T_1 ? 5'h17 : _GEN_505; // @[\\src\\main\\scala\\BlockLogic.scala 33:23 99:21]
  wire  _GEN_559 = 3'h2 == _T_1 ? 1'h0 : 3'h3 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_560 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_481); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_561 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_482); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_562 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_483); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_563 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_484); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_564 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_485); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_565 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_486); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_566 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_487); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_567 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_488); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire  _GEN_568 = 3'h2 == _T_1 ? 1'h0 : _GEN_506; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_569 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_507); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_570 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_508); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_571 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_509); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_572 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_510); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_573 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_511); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_574 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_512); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_575 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_513); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_576 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_514); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire  _GEN_577 = 3'h2 == _T_1 ? 1'h0 : _GEN_515; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_578 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_516); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_579 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_517); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_580 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_518); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_582 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_520); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_583 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_521); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_584 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_522); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_585 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_523); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire  _GEN_586 = 3'h2 == _T_1 ? 1'h0 : _GEN_524; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_587 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_525); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_588 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_526); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_589 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_527); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_590 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_528); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_591 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_529); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_592 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_530); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_593 = 3'h2 == _T_1 ? $signed(16'sh0) : $signed(_GEN_531); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_594 = 3'h2 == _T_1 ? $signed(15'sh0) : $signed(_GEN_532); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_596 = 3'h1 == _T_1 ? $signed(_GEN_26) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_597 = 3'h1 == _T_1 ? $signed(_GEN_27) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [14:0] _GEN_599 = 3'h1 == _T_1 ? $signed(_GEN_4) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_600 = 3'h1 == _T_1 ? $signed(_GEN_30) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_602 = 3'h1 == _T_1 ? $signed(_GEN_32) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_603 = 3'h1 == _T_1 ? $signed(_GEN_33) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [3:0] _GEN_604 = 3'h1 == _T_1 ? $signed(_GEN_34) : $signed(_GEN_542); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_605 = 3'h1 == _T_1 ? $signed(_GEN_34) : $signed(_GEN_543); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_606 = 3'h1 == _T_1 ? $signed(_GEN_36) : $signed(_GEN_544); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_607 = 3'h1 == _T_1 ? $signed(_GEN_37) : $signed(_GEN_545); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_608 = 3'h1 == _T_1 ? $signed(_GEN_19) : $signed(_GEN_546); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_609 = 3'h1 == _T_1 ? $signed(4'sh2) : $signed(_GEN_547); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_610 = 3'h1 == _T_1 ? $signed(4'sh2) : $signed(_GEN_548); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_611 = 3'h1 == _T_1 ? $signed(4'sh3) : $signed(_GEN_549); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_612 = 3'h1 == _T_1 ? $signed(_GEN_37) : $signed(_GEN_550); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_613 = 3'h1 == _T_1 ? $signed(_GEN_37) : $signed(_GEN_551); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_614 = 3'h1 == _T_1 ? $signed(_GEN_44) : $signed(_GEN_552); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_615 = 3'h1 == _T_1 ? $signed(_GEN_34) : $signed(_GEN_553); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_616 = 3'h1 == _T_1 ? $signed(_GEN_11) : $signed(_GEN_554); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_617 = 3'h1 == _T_1 ? $signed(4'sh2) : $signed(_GEN_555); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_618 = 3'h1 == _T_1 ? $signed(4'sh2) : $signed(_GEN_556); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [3:0] _GEN_619 = 3'h1 == _T_1 ? $signed(4'sh3) : $signed(_GEN_557); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  wire [4:0] _GEN_620 = 3'h1 == _T_1 ? 5'h16 : _GEN_558; // @[\\src\\main\\scala\\BlockLogic.scala 33:23 86:21]
  wire  _GEN_621 = 3'h1 == _T_1 ? 1'h0 : 3'h2 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_622 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_534); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_623 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_535); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [14:0] _GEN_625 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_537); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_626 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_538); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire  _GEN_630 = 3'h1 == _T_1 ? 1'h0 : _GEN_559; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_631 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_560); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_632 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_561); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_633 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_562); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_634 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_563); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_635 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_564); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_636 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_565); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_637 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_566); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_638 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_567); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire  _GEN_639 = 3'h1 == _T_1 ? 1'h0 : _GEN_568; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_640 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_569); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_641 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_570); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_642 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_571); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_643 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_572); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_644 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_573); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_645 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_574); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_646 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_575); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_647 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_576); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire  _GEN_648 = 3'h1 == _T_1 ? 1'h0 : _GEN_577; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_649 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_578); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_650 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_579); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_651 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_580); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_653 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_582); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_654 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_583); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_655 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_584); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_656 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_585); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire  _GEN_657 = 3'h1 == _T_1 ? 1'h0 : _GEN_586; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  wire [15:0] _GEN_658 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_587); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_659 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_588); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_660 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_589); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_661 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_590); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_662 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_591); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_663 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_592); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_664 = 3'h1 == _T_1 ? $signed(16'sh0) : $signed(_GEN_593); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_665 = 3'h1 == _T_1 ? $signed(15'sh0) : $signed(_GEN_594); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_667 = 3'h0 == _T_1 ? $signed(_GEN_1) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_668 = 3'h0 == _T_1 ? $signed(_GEN_2) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [14:0] _GEN_670 = 3'h0 == _T_1 ? $signed(_GEN_4) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_671 = 3'h0 == _T_1 ? $signed(_GEN_5) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_673 = 3'h0 == _T_1 ? $signed(_GEN_7) : $signed(16'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_674 = 3'h0 == _T_1 ? $signed(_GEN_8) : $signed(15'sh0); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_693 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_596); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_694 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_597); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [14:0] _GEN_696 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_599); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_697 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_600); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_699 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_602); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_700 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_603); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_702 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_622); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_703 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_623); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [14:0] _GEN_705 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_625); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_706 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_626); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_711 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_631); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_712 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_632); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_713 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_633); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_714 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_634); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_715 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_635); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_716 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_636); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_717 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_637); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_718 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_638); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_720 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_640); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_721 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_641); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_722 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_642); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_723 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_643); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_724 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_644); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_725 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_645); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_726 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_646); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_727 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_647); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_729 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_649); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_730 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_650); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_731 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_651); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [15:0] _GEN_733 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_653); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_734 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_654); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_735 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_655); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_736 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_656); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_738 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_658); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_739 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_659); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_740 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_660); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_741 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_661); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_742 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_662); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_743 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_663); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  wire [15:0] _GEN_744 = 3'h0 == _T_1 ? $signed(16'sh0) : $signed(_GEN_664); // @[\\src\\main\\scala\\BlockLogic.scala 20:22 33:23]
  wire [14:0] _GEN_745 = 3'h0 == _T_1 ? $signed(15'sh0) : $signed(_GEN_665); // @[\\src\\main\\scala\\BlockLogic.scala 21:22 33:23]
  assign io_spriteXPosition_0 = _GEN_667[10:0];
  assign io_spriteXPosition_1 = _GEN_667[10:0];
  assign io_spriteXPosition_2 = _GEN_671[10:0];
  assign io_spriteXPosition_3 = _GEN_673[10:0];
  assign io_spriteXPosition_4 = _GEN_693[10:0];
  assign io_spriteXPosition_5 = _GEN_693[10:0];
  assign io_spriteXPosition_6 = _GEN_697[10:0];
  assign io_spriteXPosition_7 = _GEN_699[10:0];
  assign io_spriteXPosition_8 = _GEN_702[10:0];
  assign io_spriteXPosition_9 = _GEN_702[10:0];
  assign io_spriteXPosition_10 = _GEN_706[10:0];
  assign io_spriteXPosition_11 = _GEN_706[10:0];
  assign io_spriteXPosition_12 = _GEN_711[10:0];
  assign io_spriteXPosition_13 = _GEN_713[10:0];
  assign io_spriteXPosition_14 = _GEN_715[10:0];
  assign io_spriteXPosition_15 = _GEN_717[10:0];
  assign io_spriteXPosition_16 = _GEN_720[10:0];
  assign io_spriteXPosition_17 = _GEN_722[10:0];
  assign io_spriteXPosition_18 = _GEN_724[10:0];
  assign io_spriteXPosition_19 = _GEN_726[10:0];
  assign io_spriteXPosition_20 = _GEN_729[10:0];
  assign io_spriteXPosition_21 = _GEN_731[10:0];
  assign io_spriteXPosition_22 = _GEN_733[10:0];
  assign io_spriteXPosition_23 = _GEN_735[10:0];
  assign io_spriteXPosition_24 = _GEN_738[10:0];
  assign io_spriteXPosition_25 = _GEN_740[10:0];
  assign io_spriteXPosition_26 = _GEN_742[10:0];
  assign io_spriteXPosition_27 = _GEN_744[10:0];
  assign io_spriteYPosition_0 = _GEN_668[9:0];
  assign io_spriteYPosition_1 = _GEN_670[9:0];
  assign io_spriteYPosition_2 = _GEN_670[9:0];
  assign io_spriteYPosition_3 = _GEN_674[9:0];
  assign io_spriteYPosition_4 = _GEN_694[9:0];
  assign io_spriteYPosition_5 = _GEN_696[9:0];
  assign io_spriteYPosition_6 = _GEN_696[9:0];
  assign io_spriteYPosition_7 = _GEN_700[9:0];
  assign io_spriteYPosition_8 = _GEN_703[9:0];
  assign io_spriteYPosition_9 = _GEN_705[9:0];
  assign io_spriteYPosition_10 = _GEN_703[9:0];
  assign io_spriteYPosition_11 = _GEN_705[9:0];
  assign io_spriteYPosition_12 = _GEN_712[9:0];
  assign io_spriteYPosition_13 = _GEN_714[9:0];
  assign io_spriteYPosition_14 = _GEN_716[9:0];
  assign io_spriteYPosition_15 = _GEN_718[9:0];
  assign io_spriteYPosition_16 = _GEN_721[9:0];
  assign io_spriteYPosition_17 = _GEN_723[9:0];
  assign io_spriteYPosition_18 = _GEN_725[9:0];
  assign io_spriteYPosition_19 = _GEN_727[9:0];
  assign io_spriteYPosition_20 = _GEN_730[9:0];
  assign io_spriteYPosition_21 = _GEN_730[9:0];
  assign io_spriteYPosition_22 = _GEN_734[9:0];
  assign io_spriteYPosition_23 = _GEN_736[9:0];
  assign io_spriteYPosition_24 = _GEN_739[9:0];
  assign io_spriteYPosition_25 = _GEN_741[9:0];
  assign io_spriteYPosition_26 = _GEN_743[9:0];
  assign io_spriteYPosition_27 = _GEN_745[9:0];
  assign io_spriteVisible_0 = 3'h0 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_spriteVisible_1 = 3'h0 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_spriteVisible_2 = 3'h0 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_spriteVisible_3 = 3'h0 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_spriteVisible_4 = 3'h0 == _T_1 ? 1'h0 : 3'h1 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_5 = 3'h0 == _T_1 ? 1'h0 : 3'h1 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_6 = 3'h0 == _T_1 ? 1'h0 : 3'h1 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_7 = 3'h0 == _T_1 ? 1'h0 : 3'h1 == _T_1; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_8 = 3'h0 == _T_1 ? 1'h0 : _GEN_621; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_9 = 3'h0 == _T_1 ? 1'h0 : _GEN_621; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_10 = 3'h0 == _T_1 ? 1'h0 : _GEN_621; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_11 = 3'h0 == _T_1 ? 1'h0 : _GEN_621; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_12 = 3'h0 == _T_1 ? 1'h0 : _GEN_630; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_13 = 3'h0 == _T_1 ? 1'h0 : _GEN_630; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_14 = 3'h0 == _T_1 ? 1'h0 : _GEN_630; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_15 = 3'h0 == _T_1 ? 1'h0 : _GEN_630; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_16 = 3'h0 == _T_1 ? 1'h0 : _GEN_639; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_17 = 3'h0 == _T_1 ? 1'h0 : _GEN_639; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_18 = 3'h0 == _T_1 ? 1'h0 : _GEN_639; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_19 = 3'h0 == _T_1 ? 1'h0 : _GEN_639; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_20 = 3'h0 == _T_1 ? 1'h0 : _GEN_648; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_21 = 3'h0 == _T_1 ? 1'h0 : _GEN_648; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_22 = 3'h0 == _T_1 ? 1'h0 : _GEN_648; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_23 = 3'h0 == _T_1 ? 1'h0 : _GEN_648; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_24 = 3'h0 == _T_1 ? 1'h0 : _GEN_657; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_25 = 3'h0 == _T_1 ? 1'h0 : _GEN_657; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_26 = 3'h0 == _T_1 ? 1'h0 : _GEN_657; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_spriteVisible_27 = 3'h0 == _T_1 ? 1'h0 : _GEN_657; // @[\\src\\main\\scala\\BlockLogic.scala 22:20 33:23]
  assign io_activeOffsetX_0 = 3'h0 == _T_1 ? $signed(4'sh2) : $signed(_GEN_604); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_activeOffsetX_1 = 3'h0 == _T_1 ? $signed(4'sh2) : $signed(_GEN_605); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_activeOffsetX_2 = 3'h0 == _T_1 ? $signed(_GEN_11) : $signed(_GEN_606); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_activeOffsetX_3 = 3'h0 == _T_1 ? $signed(4'sh3) : $signed(_GEN_607); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_activeOffsetY_0 = 3'h0 == _T_1 ? $signed(4'sh1) : $signed(_GEN_608); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_activeOffsetY_1 = 3'h0 == _T_1 ? $signed(4'sh2) : $signed(_GEN_609); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_activeOffsetY_2 = 3'h0 == _T_1 ? $signed(4'sh2) : $signed(_GEN_610); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_activeOffsetY_3 = 3'h0 == _T_1 ? $signed(_GEN_11) : $signed(_GEN_611); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_nextOffsetX_0 = 3'h0 == _T_1 ? $signed(4'sh2) : $signed(_GEN_612); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_nextOffsetX_1 = 3'h0 == _T_1 ? $signed(4'sh2) : $signed(_GEN_613); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_nextOffsetX_2 = 3'h0 == _T_1 ? $signed(_GEN_19) : $signed(_GEN_614); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_nextOffsetX_3 = 3'h0 == _T_1 ? $signed(4'sh3) : $signed(_GEN_615); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_nextOffsetY_0 = 3'h0 == _T_1 ? $signed(4'sh1) : $signed(_GEN_616); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_nextOffsetY_1 = 3'h0 == _T_1 ? $signed(4'sh2) : $signed(_GEN_617); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_nextOffsetY_2 = 3'h0 == _T_1 ? $signed(4'sh2) : $signed(_GEN_618); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_nextOffsetY_3 = 3'h0 == _T_1 ? $signed(_GEN_19) : $signed(_GEN_619); // @[\\src\\main\\scala\\BlockLogic.scala 33:23]
  assign io_tileNumber = 3'h0 == _T_1 ? 5'h15 : _GEN_620; // @[\\src\\main\\scala\\BlockLogic.scala 33:23 59:21]
endmodule
module GameLogic(
  input         clock,
  input         reset,
  input         io_btnU, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  input         io_btnL, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  input         io_btnR, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  input         io_btnD, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  input         io_sw_7, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_led_0, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_led_1, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_led_2, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_led_3, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_0, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_1, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_2, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_3, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_4, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_5, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_6, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_7, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_8, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_9, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_10, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_11, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_12, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_13, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_14, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_15, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_16, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_17, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_18, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_19, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_20, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_21, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_22, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_23, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_24, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_25, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_26, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_spriteXPosition_27, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_0, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_1, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_2, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_3, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_4, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_5, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_6, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_7, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_8, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_9, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_10, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_11, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_12, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_13, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_14, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_15, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_16, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_17, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_18, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_19, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_20, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_21, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_22, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_23, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_24, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_25, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_26, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_spriteYPosition_27, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_0, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_1, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_2, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_3, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_4, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_5, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_6, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_7, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_8, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_9, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_10, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_11, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_12, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_13, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_14, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_15, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_16, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_17, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_18, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_19, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_20, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_21, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_22, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_23, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_24, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_25, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_26, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_spriteVisible_27, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [9:0]  io_viewBoxX, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [8:0]  io_viewBoxY, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [4:0]  io_backBufferWriteData, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output [10:0] io_backBufferWriteAddress, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_backBufferWriteEnable, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  input         io_newFrame, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_frameUpdateDone, // @[\\src\\main\\scala\\GameLogic.scala 13:14]
  output        io_startTune_0 // @[\\src\\main\\scala\\GameLogic.scala 13:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] fallDetector_io_grid_0; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_1; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_2; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_3; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_4; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_5; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_6; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_7; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_8; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_9; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_10; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_11; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_12; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_13; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_14; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_15; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_16; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_17; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_18; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_19; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_20; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_21; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_22; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_23; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_24; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_25; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_26; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_27; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_28; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_29; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_30; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_31; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_32; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_33; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_34; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_35; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_36; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_37; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_38; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_39; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_40; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_41; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_42; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_43; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_44; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_45; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_46; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_47; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_48; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_49; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_50; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_51; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_52; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_53; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_54; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_55; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_56; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_57; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_58; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_59; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_60; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_61; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_62; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_63; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_64; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_65; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_66; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_67; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_68; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_69; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_70; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_71; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_72; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_73; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_74; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_75; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_76; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_77; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_78; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_79; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_80; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_81; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_82; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_83; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_84; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_85; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_86; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_87; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_88; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_89; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_90; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_91; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_92; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_93; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_94; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_95; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_96; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_97; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_98; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_99; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_100; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_101; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_102; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_103; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_104; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_105; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_106; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_107; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_108; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_109; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_110; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_111; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_112; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_113; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_114; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_115; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_116; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_117; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_118; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_119; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_120; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_121; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_122; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_123; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_124; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_125; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_126; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_127; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_128; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_129; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_130; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_131; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_132; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_133; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_134; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_135; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_136; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_137; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_138; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_139; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_140; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_141; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_142; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_143; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_144; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_145; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_146; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_147; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_148; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_149; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_150; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_151; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_152; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_153; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_154; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_155; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_156; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_157; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_158; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_159; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_160; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_161; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_162; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_163; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_164; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_165; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_166; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_167; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_168; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_169; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_170; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_171; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_172; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_173; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_174; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_175; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_176; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_177; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_178; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_179; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_180; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_181; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_182; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_183; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_184; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_185; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_186; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_187; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_188; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_189; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_190; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_191; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_192; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_193; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_194; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_195; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_196; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_197; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_198; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_199; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_200; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_201; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_202; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_203; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_204; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_205; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_206; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_207; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_208; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_209; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_210; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_211; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_212; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_213; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_214; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_215; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_216; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_217; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_218; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_219; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_220; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_221; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_222; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_223; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_224; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_225; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_226; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_227; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_228; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_229; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_230; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_231; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_232; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_233; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_234; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_235; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_236; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_237; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_238; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_239; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_240; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_241; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_242; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_243; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_244; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_245; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_246; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_247; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_248; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_249; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_250; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_251; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_252; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_253; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_254; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_255; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_256; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_257; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_258; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_259; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_260; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_261; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_262; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_263; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_264; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_265; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_266; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_267; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_268; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_269; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_270; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_271; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_272; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_273; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_274; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_275; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_276; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_277; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_278; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_279; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_280; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_281; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_282; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_283; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_284; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_285; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_286; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_287; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_288; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_289; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_290; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_291; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_292; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_293; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_294; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_295; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_296; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_297; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_298; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] fallDetector_io_grid_299; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [10:0] fallDetector_io_xPos; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [9:0] fallDetector_io_yPos; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [3:0] fallDetector_io_xOffsets_0; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [3:0] fallDetector_io_xOffsets_1; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [3:0] fallDetector_io_xOffsets_2; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [3:0] fallDetector_io_xOffsets_3; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [3:0] fallDetector_io_yOffsets_0; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [3:0] fallDetector_io_yOffsets_1; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [3:0] fallDetector_io_yOffsets_2; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [3:0] fallDetector_io_yOffsets_3; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire  fallDetector_io_isCollision; // @[\\src\\main\\scala\\GameLogic.scala 106:28]
  wire [2:0] movementDetector_io_grid_0; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_1; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_2; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_3; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_4; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_5; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_6; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_7; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_8; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_9; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_10; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_11; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_12; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_13; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_14; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_15; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_16; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_17; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_18; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_19; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_20; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_21; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_22; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_23; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_24; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_25; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_26; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_27; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_28; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_29; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_30; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_31; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_32; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_33; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_34; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_35; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_36; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_37; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_38; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_39; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_40; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_41; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_42; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_43; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_44; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_45; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_46; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_47; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_48; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_49; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_50; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_51; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_52; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_53; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_54; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_55; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_56; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_57; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_58; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_59; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_60; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_61; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_62; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_63; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_64; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_65; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_66; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_67; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_68; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_69; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_70; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_71; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_72; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_73; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_74; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_75; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_76; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_77; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_78; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_79; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_80; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_81; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_82; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_83; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_84; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_85; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_86; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_87; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_88; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_89; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_90; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_91; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_92; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_93; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_94; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_95; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_96; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_97; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_98; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_99; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_100; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_101; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_102; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_103; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_104; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_105; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_106; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_107; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_108; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_109; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_110; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_111; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_112; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_113; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_114; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_115; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_116; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_117; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_118; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_119; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_120; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_121; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_122; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_123; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_124; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_125; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_126; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_127; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_128; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_129; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_130; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_131; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_132; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_133; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_134; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_135; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_136; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_137; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_138; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_139; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_140; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_141; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_142; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_143; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_144; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_145; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_146; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_147; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_148; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_149; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_150; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_151; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_152; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_153; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_154; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_155; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_156; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_157; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_158; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_159; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_160; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_161; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_162; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_163; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_164; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_165; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_166; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_167; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_168; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_169; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_170; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_171; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_172; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_173; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_174; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_175; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_176; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_177; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_178; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_179; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_180; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_181; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_182; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_183; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_184; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_185; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_186; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_187; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_188; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_189; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_190; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_191; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_192; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_193; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_194; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_195; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_196; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_197; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_198; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_199; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_200; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_201; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_202; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_203; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_204; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_205; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_206; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_207; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_208; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_209; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_210; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_211; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_212; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_213; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_214; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_215; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_216; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_217; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_218; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_219; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_220; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_221; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_222; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_223; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_224; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_225; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_226; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_227; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_228; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_229; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_230; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_231; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_232; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_233; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_234; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_235; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_236; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_237; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_238; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_239; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_240; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_241; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_242; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_243; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_244; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_245; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_246; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_247; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_248; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_249; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_250; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_251; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_252; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_253; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_254; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_255; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_256; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_257; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_258; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_259; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_260; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_261; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_262; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_263; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_264; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_265; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_266; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_267; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_268; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_269; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_270; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_271; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_272; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_273; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_274; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_275; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_276; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_277; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_278; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_279; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_280; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_281; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_282; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_283; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_284; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_285; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_286; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_287; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_288; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_289; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_290; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_291; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_292; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_293; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_294; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_295; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_296; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_297; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_298; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [2:0] movementDetector_io_grid_299; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [10:0] movementDetector_io_xPos; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [9:0] movementDetector_io_yPos; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [3:0] movementDetector_io_xOffsets_0; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [3:0] movementDetector_io_xOffsets_1; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [3:0] movementDetector_io_xOffsets_2; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [3:0] movementDetector_io_xOffsets_3; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [3:0] movementDetector_io_yOffsets_0; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [3:0] movementDetector_io_yOffsets_1; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [3:0] movementDetector_io_yOffsets_2; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [3:0] movementDetector_io_yOffsets_3; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire  movementDetector_io_isCollision; // @[\\src\\main\\scala\\GameLogic.scala 112:32]
  wire [10:0] posToIndex_io_xPos; // @[\\src\\main\\scala\\GameLogic.scala 120:26]
  wire [9:0] posToIndex_io_yPos; // @[\\src\\main\\scala\\GameLogic.scala 120:26]
  wire [10:0] posToIndex_io_index; // @[\\src\\main\\scala\\GameLogic.scala 120:26]
  wire [10:0] posToGridIndex_io_xPos; // @[\\src\\main\\scala\\GameLogic.scala 123:30]
  wire [9:0] posToGridIndex_io_yPos; // @[\\src\\main\\scala\\GameLogic.scala 123:30]
  wire [8:0] posToGridIndex_io_index; // @[\\src\\main\\scala\\GameLogic.scala 123:30]
  wire  gameScreen_clock; // @[\\src\\main\\scala\\GameLogic.scala 151:26]
  wire  gameScreen_reset; // @[\\src\\main\\scala\\GameLogic.scala 151:26]
  wire  gameScreen_io_sw; // @[\\src\\main\\scala\\GameLogic.scala 151:26]
  wire [9:0] gameScreen_io_viewBoxX; // @[\\src\\main\\scala\\GameLogic.scala 151:26]
  wire [8:0] gameScreen_io_viewBoxY; // @[\\src\\main\\scala\\GameLogic.scala 151:26]
  wire  gameScreen_io_staticScreen; // @[\\src\\main\\scala\\GameLogic.scala 151:26]
  wire  blockType_prng_clock; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  blockType_prng_reset; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  blockType_prng_io_increment; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  blockType_prng_io_out_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  blockType_prng_io_out_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  blockType_prng_io_out_2; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  rnd_prng_clock; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  rnd_prng_reset; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  rnd_prng_io_increment; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  rnd_prng_io_out_0; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  rnd_prng_io_out_1; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire  rnd_prng_io_out_2; // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
  wire [1:0] blockLogic_io_rotation; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_xPos; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_yPos; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [2:0] blockLogic_io_sel; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_0; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_1; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_2; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_4; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_5; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_6; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_15; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [10:0] blockLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_0; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_1; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_2; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_4; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_5; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_6; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_15; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [9:0] blockLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_0; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_1; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_2; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire  blockLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_activeOffsetX_0; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_activeOffsetX_1; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_activeOffsetX_2; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_activeOffsetX_3; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_activeOffsetY_0; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_activeOffsetY_1; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_activeOffsetY_2; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_activeOffsetY_3; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_nextOffsetX_0; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_nextOffsetX_1; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_nextOffsetX_2; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_nextOffsetX_3; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_nextOffsetY_0; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_nextOffsetY_1; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_nextOffsetY_2; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [3:0] blockLogic_io_nextOffsetY_3; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  wire [4:0] blockLogic_io_tileNumber; // @[\\src\\main\\scala\\GameLogic.scala 167:26]
  reg [1:0] currentTask; // @[\\src\\main\\scala\\GameLogic.scala 80:28]
  reg [1:0] writingCount; // @[\\src\\main\\scala\\GameLogic.scala 81:29]
  reg [3:0] currentBlock; // @[\\src\\main\\scala\\GameLogic.scala 84:29]
  reg [1:0] grid_0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_1; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_2; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_3; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_4; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_5; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_6; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_7; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_8; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_9; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_10; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_11; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_12; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_13; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_14; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_15; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_16; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_17; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_18; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_19; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_20; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_21; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_22; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_23; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_24; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_25; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_26; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_27; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_28; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_29; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_30; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_31; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_32; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_33; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_34; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_35; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_36; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_37; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_38; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_39; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_40; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_41; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_42; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_43; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_44; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_45; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_46; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_47; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_48; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_49; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_50; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_51; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_52; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_53; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_54; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_55; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_56; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_57; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_58; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_59; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_60; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_61; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_62; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_63; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_64; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_65; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_66; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_67; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_68; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_69; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_70; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_71; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_72; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_73; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_74; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_75; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_76; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_77; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_78; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_79; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_80; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_81; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_82; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_83; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_84; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_85; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_86; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_87; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_88; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_89; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_90; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_91; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_92; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_93; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_94; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_95; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_96; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_97; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_98; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_99; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_100; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_101; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_102; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_103; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_104; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_105; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_106; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_107; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_108; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_109; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_110; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_111; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_112; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_113; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_114; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_115; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_116; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_117; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_118; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_119; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_120; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_121; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_122; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_123; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_124; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_125; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_126; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_127; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_128; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_129; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_130; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_131; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_132; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_133; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_134; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_135; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_136; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_137; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_138; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_139; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_140; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_141; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_142; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_143; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_144; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_145; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_146; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_147; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_148; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_149; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_150; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_151; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_152; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_153; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_154; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_155; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_156; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_157; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_158; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_159; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_160; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_161; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_162; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_163; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_164; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_165; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_166; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_167; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_168; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_169; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_170; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_171; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_172; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_173; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_174; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_175; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_176; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_177; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_178; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_179; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_180; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_181; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_182; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_183; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_184; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_185; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_186; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_187; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_188; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_189; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_190; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_191; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_192; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_193; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_194; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_195; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_196; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_197; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_198; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_199; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_200; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_201; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_202; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_203; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_204; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_205; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_206; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_207; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_208; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_209; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_210; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_211; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_212; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_213; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_214; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_215; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_216; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_217; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_218; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_219; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_220; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_221; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_222; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_223; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_224; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_225; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_226; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_227; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_228; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_229; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_230; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_231; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_232; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_233; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_234; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_235; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_236; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_237; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_238; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_239; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_240; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_241; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_242; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_243; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_244; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_245; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_246; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_247; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_248; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_249; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_250; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_251; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_252; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_253; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_254; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_255; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_256; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_257; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_258; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_259; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_260; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_261; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_262; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_263; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_264; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_265; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_266; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_267; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_268; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_269; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_270; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_271; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_272; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_273; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_274; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_275; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_276; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_277; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_278; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_279; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_280; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_281; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_282; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_283; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_284; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_285; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_286; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_287; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_288; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_289; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_290; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_291; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_292; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_293; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_294; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_295; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_296; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_297; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_298; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [1:0] grid_299; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
  reg [10:0] blockXReg; // @[\\src\\main\\scala\\GameLogic.scala 102:26]
  reg [9:0] blockYReg; // @[\\src\\main\\scala\\GameLogic.scala 103:26]
  reg [1:0] stateReg; // @[\\src\\main\\scala\\GameLogic.scala 137:25]
  reg [6:0] moveCnt; // @[\\src\\main\\scala\\GameLogic.scala 142:24]
  reg [1:0] rotation; // @[\\src\\main\\scala\\GameLogic.scala 147:25]
  reg  upRelease; // @[\\src\\main\\scala\\GameLogic.scala 149:26]
  wire [2:0] _blockType_T = {blockType_prng_io_out_2,blockType_prng_io_out_1,blockType_prng_io_out_0}; // @[src/main/scala/chisel3/util/random/PRNG.scala 95:17]
  reg [2:0] blockType; // @[\\src\\main\\scala\\GameLogic.scala 157:26]
  wire [2:0] rnd = {rnd_prng_io_out_2,rnd_prng_io_out_1,rnd_prng_io_out_0}; // @[src/main/scala/chisel3/util/random/PRNG.scala 95:17]
  reg  newPiece; // @[\\src\\main\\scala\\GameLogic.scala 165:25]
  reg [6:0] speedThreshold; // @[\\src\\main\\scala\\GameLogic.scala 178:31]
  wire  _T_4 = 2'h1 == currentTask; // @[\\src\\main\\scala\\GameLogic.scala 196:27]
  wire [3:0] _GEN_2 = blockLogic_io_activeOffsetX_0; // @[\\src\\main\\scala\\GameLogic.scala 199:{47,47}]
  wire [3:0] _GEN_3 = 2'h1 == writingCount ? $signed(blockLogic_io_activeOffsetX_1) : $signed(_GEN_2); // @[\\src\\main\\scala\\GameLogic.scala 199:{47,47}]
  wire [3:0] _GEN_4 = 2'h2 == writingCount ? $signed(blockLogic_io_activeOffsetX_2) : $signed(_GEN_3); // @[\\src\\main\\scala\\GameLogic.scala 199:{47,47}]
  wire [3:0] _GEN_5 = 2'h3 == writingCount ? $signed(blockLogic_io_activeOffsetX_3) : $signed(_GEN_4); // @[\\src\\main\\scala\\GameLogic.scala 199:{47,47}]
  wire [10:0] _GEN_3492 = {{7{_GEN_5[3]}},_GEN_5}; // @[\\src\\main\\scala\\GameLogic.scala 199:47]
  wire [10:0] _posToGridIndex_io_xPos_T_2 = $signed(blockXReg) + $signed(_GEN_3492); // @[\\src\\main\\scala\\GameLogic.scala 199:47]
  wire [3:0] _GEN_6 = blockLogic_io_activeOffsetY_0; // @[\\src\\main\\scala\\GameLogic.scala 200:{47,47}]
  wire [3:0] _GEN_7 = 2'h1 == writingCount ? $signed(blockLogic_io_activeOffsetY_1) : $signed(_GEN_6); // @[\\src\\main\\scala\\GameLogic.scala 200:{47,47}]
  wire [3:0] _GEN_8 = 2'h2 == writingCount ? $signed(blockLogic_io_activeOffsetY_2) : $signed(_GEN_7); // @[\\src\\main\\scala\\GameLogic.scala 200:{47,47}]
  wire [3:0] _GEN_9 = 2'h3 == writingCount ? $signed(blockLogic_io_activeOffsetY_3) : $signed(_GEN_8); // @[\\src\\main\\scala\\GameLogic.scala 200:{47,47}]
  wire [9:0] _GEN_3493 = {{6{_GEN_9[3]}},_GEN_9}; // @[\\src\\main\\scala\\GameLogic.scala 200:47]
  wire [9:0] _posToGridIndex_io_yPos_T_2 = $signed(blockYReg) + $signed(_GEN_3493); // @[\\src\\main\\scala\\GameLogic.scala 200:47]
  wire [4:0] _grid_T_1 = 5'h14 - blockLogic_io_tileNumber; // @[\\src\\main\\scala\\GameLogic.scala 203:49]
  wire [1:0] _GEN_10 = 9'h0 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_11 = 9'h1 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_12 = 9'h2 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_13 = 9'h3 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_14 = 9'h4 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_15 = 9'h5 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_16 = 9'h6 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_17 = 9'h7 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_18 = 9'h8 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_19 = 9'h9 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_20 = 9'ha == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_21 = 9'hb == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_22 = 9'hc == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_23 = 9'hd == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_24 = 9'he == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_25 = 9'hf == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_26 = 9'h10 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_27 = 9'h11 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_28 = 9'h12 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_29 = 9'h13 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_30 = 9'h14 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_31 = 9'h15 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_32 = 9'h16 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_33 = 9'h17 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_34 = 9'h18 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 95:13]
  wire [1:0] _GEN_35 = 9'h19 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_25; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_36 = 9'h1a == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_26; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_37 = 9'h1b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_27; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_38 = 9'h1c == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_28; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_39 = 9'h1d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_29; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_40 = 9'h1e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_30; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_41 = 9'h1f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_31; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_42 = 9'h20 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_32; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_43 = 9'h21 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_33; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_44 = 9'h22 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_34; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_45 = 9'h23 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_35; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_46 = 9'h24 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_36; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_47 = 9'h25 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_37; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_48 = 9'h26 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_38; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_49 = 9'h27 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_39; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_50 = 9'h28 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_40; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_51 = 9'h29 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_41; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_52 = 9'h2a == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_42; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_53 = 9'h2b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_43; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_54 = 9'h2c == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_44; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_55 = 9'h2d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_45; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_56 = 9'h2e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_46; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_57 = 9'h2f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_47; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_58 = 9'h30 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_48; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_59 = 9'h31 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_60 = 9'h32 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_50; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_61 = 9'h33 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_51; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_62 = 9'h34 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_52; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_63 = 9'h35 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_53; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_64 = 9'h36 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_54; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_65 = 9'h37 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_55; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_66 = 9'h38 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_56; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_67 = 9'h39 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_57; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_68 = 9'h3a == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_58; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_69 = 9'h3b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_59; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_70 = 9'h3c == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_60; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_71 = 9'h3d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_61; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_72 = 9'h3e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_62; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_73 = 9'h3f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_63; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_74 = 9'h40 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_64; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_75 = 9'h41 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_65; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_76 = 9'h42 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_66; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_77 = 9'h43 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_67; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_78 = 9'h44 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_68; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_79 = 9'h45 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_69; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_80 = 9'h46 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_70; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_81 = 9'h47 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_71; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_82 = 9'h48 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_72; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_83 = 9'h49 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_73; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_84 = 9'h4a == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_85 = 9'h4b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_75; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_86 = 9'h4c == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_76; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_87 = 9'h4d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_77; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_88 = 9'h4e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_78; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_89 = 9'h4f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_79; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_90 = 9'h50 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_80; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_91 = 9'h51 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_81; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_92 = 9'h52 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_82; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_93 = 9'h53 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_83; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_94 = 9'h54 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_84; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_95 = 9'h55 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_85; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_96 = 9'h56 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_86; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_97 = 9'h57 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_87; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_98 = 9'h58 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_88; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_99 = 9'h59 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_89; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_100 = 9'h5a == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_90; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_101 = 9'h5b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_91; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_102 = 9'h5c == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_92; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_103 = 9'h5d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_93; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_104 = 9'h5e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_94; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_105 = 9'h5f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_95; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_106 = 9'h60 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_96; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_107 = 9'h61 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_97; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_108 = 9'h62 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_98; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_109 = 9'h63 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_110 = 9'h64 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_100; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_111 = 9'h65 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_101; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_112 = 9'h66 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_102; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_113 = 9'h67 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_103; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_114 = 9'h68 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_104; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_115 = 9'h69 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_105; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_116 = 9'h6a == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_106; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_117 = 9'h6b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_107; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_118 = 9'h6c == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_108; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_119 = 9'h6d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_109; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_120 = 9'h6e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_110; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_121 = 9'h6f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_111; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_122 = 9'h70 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_112; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_123 = 9'h71 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_113; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_124 = 9'h72 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_114; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_125 = 9'h73 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_115; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_126 = 9'h74 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_116; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_127 = 9'h75 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_117; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_128 = 9'h76 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_118; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_129 = 9'h77 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_119; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_130 = 9'h78 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_120; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_131 = 9'h79 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_121; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_132 = 9'h7a == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_122; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_133 = 9'h7b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_123; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_134 = 9'h7c == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_135 = 9'h7d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_125; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_136 = 9'h7e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_126; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_137 = 9'h7f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_127; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_138 = 9'h80 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_128; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_139 = 9'h81 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_129; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_140 = 9'h82 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_130; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_141 = 9'h83 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_131; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_142 = 9'h84 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_132; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_143 = 9'h85 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_133; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_144 = 9'h86 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_134; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_145 = 9'h87 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_135; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_146 = 9'h88 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_136; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_147 = 9'h89 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_137; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_148 = 9'h8a == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_138; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_149 = 9'h8b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_139; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_150 = 9'h8c == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_140; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_151 = 9'h8d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_141; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_152 = 9'h8e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_142; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_153 = 9'h8f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_143; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_154 = 9'h90 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_144; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_155 = 9'h91 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_145; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_156 = 9'h92 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_146; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_157 = 9'h93 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_147; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_158 = 9'h94 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_148; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_159 = 9'h95 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_160 = 9'h96 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_150; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_161 = 9'h97 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_151; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_162 = 9'h98 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_152; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_163 = 9'h99 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_153; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_164 = 9'h9a == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_154; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_165 = 9'h9b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_155; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_166 = 9'h9c == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_156; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_167 = 9'h9d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_157; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_168 = 9'h9e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_158; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_169 = 9'h9f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_159; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_170 = 9'ha0 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_160; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_171 = 9'ha1 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_161; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_172 = 9'ha2 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_162; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_173 = 9'ha3 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_163; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_174 = 9'ha4 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_164; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_175 = 9'ha5 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_165; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_176 = 9'ha6 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_166; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_177 = 9'ha7 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_167; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_178 = 9'ha8 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_168; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_179 = 9'ha9 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_169; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_180 = 9'haa == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_170; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_181 = 9'hab == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_171; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_182 = 9'hac == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_172; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_183 = 9'had == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_173; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_184 = 9'hae == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_185 = 9'haf == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_175; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_186 = 9'hb0 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_176; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_187 = 9'hb1 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_177; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_188 = 9'hb2 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_178; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_189 = 9'hb3 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_179; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_190 = 9'hb4 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_180; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_191 = 9'hb5 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_181; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_192 = 9'hb6 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_182; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_193 = 9'hb7 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_183; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_194 = 9'hb8 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_184; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_195 = 9'hb9 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_185; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_196 = 9'hba == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_186; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_197 = 9'hbb == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_187; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_198 = 9'hbc == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_188; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_199 = 9'hbd == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_189; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_200 = 9'hbe == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_190; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_201 = 9'hbf == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_191; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_202 = 9'hc0 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_192; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_203 = 9'hc1 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_193; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_204 = 9'hc2 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_194; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_205 = 9'hc3 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_195; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_206 = 9'hc4 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_196; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_207 = 9'hc5 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_197; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_208 = 9'hc6 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_198; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_209 = 9'hc7 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_210 = 9'hc8 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_200; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_211 = 9'hc9 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_201; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_212 = 9'hca == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_202; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_213 = 9'hcb == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_203; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_214 = 9'hcc == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_204; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_215 = 9'hcd == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_205; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_216 = 9'hce == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_206; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_217 = 9'hcf == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_207; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_218 = 9'hd0 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_208; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_219 = 9'hd1 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_209; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_220 = 9'hd2 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_210; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_221 = 9'hd3 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_211; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_222 = 9'hd4 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_212; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_223 = 9'hd5 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_213; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_224 = 9'hd6 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_214; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_225 = 9'hd7 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_215; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_226 = 9'hd8 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_216; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_227 = 9'hd9 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_217; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_228 = 9'hda == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_218; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_229 = 9'hdb == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_219; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_230 = 9'hdc == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_220; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_231 = 9'hdd == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_221; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_232 = 9'hde == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_222; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_233 = 9'hdf == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_223; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_234 = 9'he0 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_235 = 9'he1 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_225; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_236 = 9'he2 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_226; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_237 = 9'he3 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_227; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_238 = 9'he4 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_228; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_239 = 9'he5 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_229; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_240 = 9'he6 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_230; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_241 = 9'he7 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_231; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_242 = 9'he8 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_232; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_243 = 9'he9 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_233; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_244 = 9'hea == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_234; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_245 = 9'heb == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_235; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_246 = 9'hec == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_236; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_247 = 9'hed == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_237; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_248 = 9'hee == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_238; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_249 = 9'hef == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_239; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_250 = 9'hf0 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_240; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_251 = 9'hf1 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_241; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_252 = 9'hf2 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_242; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_253 = 9'hf3 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_243; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_254 = 9'hf4 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_244; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_255 = 9'hf5 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_245; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_256 = 9'hf6 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_246; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_257 = 9'hf7 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_247; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_258 = 9'hf8 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_248; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_259 = 9'hf9 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_260 = 9'hfa == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_250; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_261 = 9'hfb == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_251; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_262 = 9'hfc == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_252; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_263 = 9'hfd == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_253; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_264 = 9'hfe == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_254; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_265 = 9'hff == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_255; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_266 = 9'h100 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_256; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_267 = 9'h101 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_257; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_268 = 9'h102 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_258; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_269 = 9'h103 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_259; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_270 = 9'h104 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_260; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_271 = 9'h105 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_261; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_272 = 9'h106 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_262; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_273 = 9'h107 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_263; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_274 = 9'h108 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_264; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_275 = 9'h109 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_265; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_276 = 9'h10a == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_266; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_277 = 9'h10b == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_267; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_278 = 9'h10c == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_268; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_279 = 9'h10d == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_269; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_280 = 9'h10e == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_270; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_281 = 9'h10f == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_271; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_282 = 9'h110 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_272; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_283 = 9'h111 == posToGridIndex_io_index ? _grid_T_1[1:0] : grid_273; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 88:21]
  wire [1:0] _GEN_284 = 9'h112 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 91:23]
  wire [1:0] _GEN_285 = 9'h113 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_286 = 9'h114 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_287 = 9'h115 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_288 = 9'h116 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_289 = 9'h117 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_290 = 9'h118 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_291 = 9'h119 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_292 = 9'h11a == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_293 = 9'h11b == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_294 = 9'h11c == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_295 = 9'h11d == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_296 = 9'h11e == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_297 = 9'h11f == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_298 = 9'h120 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_299 = 9'h121 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_300 = 9'h122 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_301 = 9'h123 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_302 = 9'h124 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_303 = 9'h125 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_304 = 9'h126 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_305 = 9'h127 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_306 = 9'h128 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_307 = 9'h129 == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_308 = 9'h12a == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _GEN_309 = 9'h12b == posToGridIndex_io_index ? _grid_T_1[1:0] : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 203:{41,41} 96:21]
  wire [1:0] _writingCount_T_1 = writingCount + 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 215:53]
  wire [1:0] _GEN_310 = writingCount == 2'h3 ? 2'h0 : _writingCount_T_1; // @[\\src\\main\\scala\\GameLogic.scala 206:38 207:26 215:37]
  wire [10:0] _GEN_311 = writingCount == 2'h3 ? $signed(-11'sh4) : $signed(blockXReg); // @[\\src\\main\\scala\\GameLogic.scala 206:38 208:23 102:26]
  wire [9:0] _GEN_312 = writingCount == 2'h3 ? $signed(10'sh8) : $signed(blockYReg); // @[\\src\\main\\scala\\GameLogic.scala 206:38 209:23 103:26]
  wire [1:0] _GEN_313 = writingCount == 2'h3 ? 2'h0 : currentTask; // @[\\src\\main\\scala\\GameLogic.scala 206:38 210:25 80:28]
  wire [1:0] _GEN_314 = writingCount == 2'h3 ? 2'h3 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 206:38 211:22 137:25]
  wire  _GEN_315 = writingCount == 2'h3 | newPiece; // @[\\src\\main\\scala\\GameLogic.scala 206:38 212:22 165:25]
  wire [1:0] _GEN_316 = writingCount == 2'h3 ? 2'h0 : rotation; // @[\\src\\main\\scala\\GameLogic.scala 206:38 213:22 147:25]
  wire [8:0] _GEN_318 = 4'h1 == currentBlock ? 9'h78 : 9'h64; // @[\\src\\main\\scala\\GameLogic.scala 225:{51,51}]
  wire [8:0] _GEN_319 = 4'h2 == currentBlock ? 9'h8c : _GEN_318; // @[\\src\\main\\scala\\GameLogic.scala 225:{51,51}]
  wire [8:0] _GEN_320 = 4'h3 == currentBlock ? 9'ha0 : _GEN_319; // @[\\src\\main\\scala\\GameLogic.scala 225:{51,51}]
  wire [8:0] _GEN_321 = 4'h4 == currentBlock ? 9'hb4 : _GEN_320; // @[\\src\\main\\scala\\GameLogic.scala 225:{51,51}]
  wire [8:0] _GEN_322 = 4'h5 == currentBlock ? 9'hc8 : _GEN_321; // @[\\src\\main\\scala\\GameLogic.scala 225:{51,51}]
  wire [8:0] _GEN_323 = 4'h6 == currentBlock ? 9'hdc : _GEN_322; // @[\\src\\main\\scala\\GameLogic.scala 225:{51,51}]
  wire [8:0] _GEN_324 = 4'h7 == currentBlock ? 9'hf0 : _GEN_323; // @[\\src\\main\\scala\\GameLogic.scala 225:{51,51}]
  wire [8:0] _GEN_325 = 4'h8 == currentBlock ? 9'h104 : _GEN_324; // @[\\src\\main\\scala\\GameLogic.scala 225:{51,51}]
  wire [8:0] _GEN_326 = 4'h9 == currentBlock ? 9'h118 : _GEN_325; // @[\\src\\main\\scala\\GameLogic.scala 225:{51,51}]
  wire [9:0] _index_T = {{1'd0}, _GEN_326}; // @[\\src\\main\\scala\\GameLogic.scala 225:51]
  wire [8:0] index = _index_T[8:0]; // @[\\src\\main\\scala\\GameLogic.scala 225:51]
  wire [8:0] _aboveValue_T_1 = index - 9'h1; // @[\\src\\main\\scala\\GameLogic.scala 227:41]
  wire [1:0] _GEN_328 = 9'h1 == index ? grid_1 : grid_0; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_329 = 9'h2 == index ? grid_2 : _GEN_328; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_330 = 9'h3 == index ? grid_3 : _GEN_329; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_331 = 9'h4 == index ? grid_4 : _GEN_330; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_332 = 9'h5 == index ? grid_5 : _GEN_331; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_333 = 9'h6 == index ? grid_6 : _GEN_332; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_334 = 9'h7 == index ? grid_7 : _GEN_333; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_335 = 9'h8 == index ? grid_8 : _GEN_334; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_336 = 9'h9 == index ? grid_9 : _GEN_335; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_337 = 9'ha == index ? grid_10 : _GEN_336; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_338 = 9'hb == index ? grid_11 : _GEN_337; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_339 = 9'hc == index ? grid_12 : _GEN_338; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_340 = 9'hd == index ? grid_13 : _GEN_339; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_341 = 9'he == index ? grid_14 : _GEN_340; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_342 = 9'hf == index ? grid_15 : _GEN_341; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_343 = 9'h10 == index ? grid_16 : _GEN_342; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_344 = 9'h11 == index ? grid_17 : _GEN_343; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_345 = 9'h12 == index ? grid_18 : _GEN_344; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_346 = 9'h13 == index ? grid_19 : _GEN_345; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_347 = 9'h14 == index ? grid_20 : _GEN_346; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_348 = 9'h15 == index ? grid_21 : _GEN_347; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_349 = 9'h16 == index ? grid_22 : _GEN_348; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_350 = 9'h17 == index ? grid_23 : _GEN_349; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_351 = 9'h18 == index ? grid_24 : _GEN_350; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_352 = 9'h19 == index ? grid_25 : _GEN_351; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_353 = 9'h1a == index ? grid_26 : _GEN_352; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_354 = 9'h1b == index ? grid_27 : _GEN_353; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_355 = 9'h1c == index ? grid_28 : _GEN_354; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_356 = 9'h1d == index ? grid_29 : _GEN_355; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_357 = 9'h1e == index ? grid_30 : _GEN_356; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_358 = 9'h1f == index ? grid_31 : _GEN_357; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_359 = 9'h20 == index ? grid_32 : _GEN_358; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_360 = 9'h21 == index ? grid_33 : _GEN_359; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_361 = 9'h22 == index ? grid_34 : _GEN_360; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_362 = 9'h23 == index ? grid_35 : _GEN_361; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_363 = 9'h24 == index ? grid_36 : _GEN_362; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_364 = 9'h25 == index ? grid_37 : _GEN_363; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_365 = 9'h26 == index ? grid_38 : _GEN_364; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_366 = 9'h27 == index ? grid_39 : _GEN_365; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_367 = 9'h28 == index ? grid_40 : _GEN_366; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_368 = 9'h29 == index ? grid_41 : _GEN_367; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_369 = 9'h2a == index ? grid_42 : _GEN_368; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_370 = 9'h2b == index ? grid_43 : _GEN_369; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_371 = 9'h2c == index ? grid_44 : _GEN_370; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_372 = 9'h2d == index ? grid_45 : _GEN_371; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_373 = 9'h2e == index ? grid_46 : _GEN_372; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_374 = 9'h2f == index ? grid_47 : _GEN_373; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_375 = 9'h30 == index ? grid_48 : _GEN_374; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_376 = 9'h31 == index ? grid_49 : _GEN_375; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_377 = 9'h32 == index ? grid_50 : _GEN_376; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_378 = 9'h33 == index ? grid_51 : _GEN_377; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_379 = 9'h34 == index ? grid_52 : _GEN_378; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_380 = 9'h35 == index ? grid_53 : _GEN_379; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_381 = 9'h36 == index ? grid_54 : _GEN_380; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_382 = 9'h37 == index ? grid_55 : _GEN_381; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_383 = 9'h38 == index ? grid_56 : _GEN_382; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_384 = 9'h39 == index ? grid_57 : _GEN_383; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_385 = 9'h3a == index ? grid_58 : _GEN_384; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_386 = 9'h3b == index ? grid_59 : _GEN_385; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_387 = 9'h3c == index ? grid_60 : _GEN_386; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_388 = 9'h3d == index ? grid_61 : _GEN_387; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_389 = 9'h3e == index ? grid_62 : _GEN_388; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_390 = 9'h3f == index ? grid_63 : _GEN_389; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_391 = 9'h40 == index ? grid_64 : _GEN_390; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_392 = 9'h41 == index ? grid_65 : _GEN_391; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_393 = 9'h42 == index ? grid_66 : _GEN_392; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_394 = 9'h43 == index ? grid_67 : _GEN_393; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_395 = 9'h44 == index ? grid_68 : _GEN_394; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_396 = 9'h45 == index ? grid_69 : _GEN_395; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_397 = 9'h46 == index ? grid_70 : _GEN_396; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_398 = 9'h47 == index ? grid_71 : _GEN_397; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_399 = 9'h48 == index ? grid_72 : _GEN_398; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_400 = 9'h49 == index ? grid_73 : _GEN_399; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_401 = 9'h4a == index ? grid_74 : _GEN_400; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_402 = 9'h4b == index ? grid_75 : _GEN_401; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_403 = 9'h4c == index ? grid_76 : _GEN_402; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_404 = 9'h4d == index ? grid_77 : _GEN_403; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_405 = 9'h4e == index ? grid_78 : _GEN_404; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_406 = 9'h4f == index ? grid_79 : _GEN_405; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_407 = 9'h50 == index ? grid_80 : _GEN_406; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_408 = 9'h51 == index ? grid_81 : _GEN_407; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_409 = 9'h52 == index ? grid_82 : _GEN_408; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_410 = 9'h53 == index ? grid_83 : _GEN_409; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_411 = 9'h54 == index ? grid_84 : _GEN_410; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_412 = 9'h55 == index ? grid_85 : _GEN_411; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_413 = 9'h56 == index ? grid_86 : _GEN_412; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_414 = 9'h57 == index ? grid_87 : _GEN_413; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_415 = 9'h58 == index ? grid_88 : _GEN_414; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_416 = 9'h59 == index ? grid_89 : _GEN_415; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_417 = 9'h5a == index ? grid_90 : _GEN_416; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_418 = 9'h5b == index ? grid_91 : _GEN_417; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_419 = 9'h5c == index ? grid_92 : _GEN_418; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_420 = 9'h5d == index ? grid_93 : _GEN_419; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_421 = 9'h5e == index ? grid_94 : _GEN_420; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_422 = 9'h5f == index ? grid_95 : _GEN_421; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_423 = 9'h60 == index ? grid_96 : _GEN_422; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_424 = 9'h61 == index ? grid_97 : _GEN_423; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_425 = 9'h62 == index ? grid_98 : _GEN_424; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_426 = 9'h63 == index ? grid_99 : _GEN_425; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_427 = 9'h64 == index ? grid_100 : _GEN_426; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_428 = 9'h65 == index ? grid_101 : _GEN_427; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_429 = 9'h66 == index ? grid_102 : _GEN_428; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_430 = 9'h67 == index ? grid_103 : _GEN_429; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_431 = 9'h68 == index ? grid_104 : _GEN_430; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_432 = 9'h69 == index ? grid_105 : _GEN_431; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_433 = 9'h6a == index ? grid_106 : _GEN_432; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_434 = 9'h6b == index ? grid_107 : _GEN_433; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_435 = 9'h6c == index ? grid_108 : _GEN_434; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_436 = 9'h6d == index ? grid_109 : _GEN_435; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_437 = 9'h6e == index ? grid_110 : _GEN_436; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_438 = 9'h6f == index ? grid_111 : _GEN_437; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_439 = 9'h70 == index ? grid_112 : _GEN_438; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_440 = 9'h71 == index ? grid_113 : _GEN_439; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_441 = 9'h72 == index ? grid_114 : _GEN_440; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_442 = 9'h73 == index ? grid_115 : _GEN_441; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_443 = 9'h74 == index ? grid_116 : _GEN_442; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_444 = 9'h75 == index ? grid_117 : _GEN_443; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_445 = 9'h76 == index ? grid_118 : _GEN_444; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_446 = 9'h77 == index ? grid_119 : _GEN_445; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_447 = 9'h78 == index ? grid_120 : _GEN_446; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_448 = 9'h79 == index ? grid_121 : _GEN_447; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_449 = 9'h7a == index ? grid_122 : _GEN_448; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_450 = 9'h7b == index ? grid_123 : _GEN_449; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_451 = 9'h7c == index ? grid_124 : _GEN_450; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_452 = 9'h7d == index ? grid_125 : _GEN_451; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_453 = 9'h7e == index ? grid_126 : _GEN_452; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_454 = 9'h7f == index ? grid_127 : _GEN_453; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_455 = 9'h80 == index ? grid_128 : _GEN_454; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_456 = 9'h81 == index ? grid_129 : _GEN_455; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_457 = 9'h82 == index ? grid_130 : _GEN_456; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_458 = 9'h83 == index ? grid_131 : _GEN_457; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_459 = 9'h84 == index ? grid_132 : _GEN_458; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_460 = 9'h85 == index ? grid_133 : _GEN_459; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_461 = 9'h86 == index ? grid_134 : _GEN_460; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_462 = 9'h87 == index ? grid_135 : _GEN_461; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_463 = 9'h88 == index ? grid_136 : _GEN_462; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_464 = 9'h89 == index ? grid_137 : _GEN_463; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_465 = 9'h8a == index ? grid_138 : _GEN_464; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_466 = 9'h8b == index ? grid_139 : _GEN_465; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_467 = 9'h8c == index ? grid_140 : _GEN_466; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_468 = 9'h8d == index ? grid_141 : _GEN_467; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_469 = 9'h8e == index ? grid_142 : _GEN_468; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_470 = 9'h8f == index ? grid_143 : _GEN_469; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_471 = 9'h90 == index ? grid_144 : _GEN_470; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_472 = 9'h91 == index ? grid_145 : _GEN_471; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_473 = 9'h92 == index ? grid_146 : _GEN_472; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_474 = 9'h93 == index ? grid_147 : _GEN_473; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_475 = 9'h94 == index ? grid_148 : _GEN_474; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_476 = 9'h95 == index ? grid_149 : _GEN_475; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_477 = 9'h96 == index ? grid_150 : _GEN_476; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_478 = 9'h97 == index ? grid_151 : _GEN_477; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_479 = 9'h98 == index ? grid_152 : _GEN_478; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_480 = 9'h99 == index ? grid_153 : _GEN_479; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_481 = 9'h9a == index ? grid_154 : _GEN_480; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_482 = 9'h9b == index ? grid_155 : _GEN_481; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_483 = 9'h9c == index ? grid_156 : _GEN_482; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_484 = 9'h9d == index ? grid_157 : _GEN_483; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_485 = 9'h9e == index ? grid_158 : _GEN_484; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_486 = 9'h9f == index ? grid_159 : _GEN_485; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_487 = 9'ha0 == index ? grid_160 : _GEN_486; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_488 = 9'ha1 == index ? grid_161 : _GEN_487; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_489 = 9'ha2 == index ? grid_162 : _GEN_488; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_490 = 9'ha3 == index ? grid_163 : _GEN_489; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_491 = 9'ha4 == index ? grid_164 : _GEN_490; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_492 = 9'ha5 == index ? grid_165 : _GEN_491; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_493 = 9'ha6 == index ? grid_166 : _GEN_492; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_494 = 9'ha7 == index ? grid_167 : _GEN_493; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_495 = 9'ha8 == index ? grid_168 : _GEN_494; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_496 = 9'ha9 == index ? grid_169 : _GEN_495; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_497 = 9'haa == index ? grid_170 : _GEN_496; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_498 = 9'hab == index ? grid_171 : _GEN_497; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_499 = 9'hac == index ? grid_172 : _GEN_498; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_500 = 9'had == index ? grid_173 : _GEN_499; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_501 = 9'hae == index ? grid_174 : _GEN_500; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_502 = 9'haf == index ? grid_175 : _GEN_501; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_503 = 9'hb0 == index ? grid_176 : _GEN_502; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_504 = 9'hb1 == index ? grid_177 : _GEN_503; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_505 = 9'hb2 == index ? grid_178 : _GEN_504; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_506 = 9'hb3 == index ? grid_179 : _GEN_505; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_507 = 9'hb4 == index ? grid_180 : _GEN_506; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_508 = 9'hb5 == index ? grid_181 : _GEN_507; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_509 = 9'hb6 == index ? grid_182 : _GEN_508; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_510 = 9'hb7 == index ? grid_183 : _GEN_509; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_511 = 9'hb8 == index ? grid_184 : _GEN_510; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_512 = 9'hb9 == index ? grid_185 : _GEN_511; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_513 = 9'hba == index ? grid_186 : _GEN_512; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_514 = 9'hbb == index ? grid_187 : _GEN_513; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_515 = 9'hbc == index ? grid_188 : _GEN_514; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_516 = 9'hbd == index ? grid_189 : _GEN_515; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_517 = 9'hbe == index ? grid_190 : _GEN_516; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_518 = 9'hbf == index ? grid_191 : _GEN_517; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_519 = 9'hc0 == index ? grid_192 : _GEN_518; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_520 = 9'hc1 == index ? grid_193 : _GEN_519; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_521 = 9'hc2 == index ? grid_194 : _GEN_520; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_522 = 9'hc3 == index ? grid_195 : _GEN_521; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_523 = 9'hc4 == index ? grid_196 : _GEN_522; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_524 = 9'hc5 == index ? grid_197 : _GEN_523; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_525 = 9'hc6 == index ? grid_198 : _GEN_524; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_526 = 9'hc7 == index ? grid_199 : _GEN_525; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_527 = 9'hc8 == index ? grid_200 : _GEN_526; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_528 = 9'hc9 == index ? grid_201 : _GEN_527; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_529 = 9'hca == index ? grid_202 : _GEN_528; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_530 = 9'hcb == index ? grid_203 : _GEN_529; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_531 = 9'hcc == index ? grid_204 : _GEN_530; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_532 = 9'hcd == index ? grid_205 : _GEN_531; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_533 = 9'hce == index ? grid_206 : _GEN_532; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_534 = 9'hcf == index ? grid_207 : _GEN_533; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_535 = 9'hd0 == index ? grid_208 : _GEN_534; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_536 = 9'hd1 == index ? grid_209 : _GEN_535; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_537 = 9'hd2 == index ? grid_210 : _GEN_536; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_538 = 9'hd3 == index ? grid_211 : _GEN_537; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_539 = 9'hd4 == index ? grid_212 : _GEN_538; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_540 = 9'hd5 == index ? grid_213 : _GEN_539; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_541 = 9'hd6 == index ? grid_214 : _GEN_540; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_542 = 9'hd7 == index ? grid_215 : _GEN_541; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_543 = 9'hd8 == index ? grid_216 : _GEN_542; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_544 = 9'hd9 == index ? grid_217 : _GEN_543; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_545 = 9'hda == index ? grid_218 : _GEN_544; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_546 = 9'hdb == index ? grid_219 : _GEN_545; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_547 = 9'hdc == index ? grid_220 : _GEN_546; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_548 = 9'hdd == index ? grid_221 : _GEN_547; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_549 = 9'hde == index ? grid_222 : _GEN_548; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_550 = 9'hdf == index ? grid_223 : _GEN_549; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_551 = 9'he0 == index ? grid_224 : _GEN_550; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_552 = 9'he1 == index ? grid_225 : _GEN_551; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_553 = 9'he2 == index ? grid_226 : _GEN_552; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_554 = 9'he3 == index ? grid_227 : _GEN_553; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_555 = 9'he4 == index ? grid_228 : _GEN_554; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_556 = 9'he5 == index ? grid_229 : _GEN_555; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_557 = 9'he6 == index ? grid_230 : _GEN_556; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_558 = 9'he7 == index ? grid_231 : _GEN_557; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_559 = 9'he8 == index ? grid_232 : _GEN_558; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_560 = 9'he9 == index ? grid_233 : _GEN_559; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_561 = 9'hea == index ? grid_234 : _GEN_560; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_562 = 9'heb == index ? grid_235 : _GEN_561; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_563 = 9'hec == index ? grid_236 : _GEN_562; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_564 = 9'hed == index ? grid_237 : _GEN_563; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_565 = 9'hee == index ? grid_238 : _GEN_564; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_566 = 9'hef == index ? grid_239 : _GEN_565; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_567 = 9'hf0 == index ? grid_240 : _GEN_566; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_568 = 9'hf1 == index ? grid_241 : _GEN_567; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_569 = 9'hf2 == index ? grid_242 : _GEN_568; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_570 = 9'hf3 == index ? grid_243 : _GEN_569; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_571 = 9'hf4 == index ? grid_244 : _GEN_570; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_572 = 9'hf5 == index ? grid_245 : _GEN_571; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_573 = 9'hf6 == index ? grid_246 : _GEN_572; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_574 = 9'hf7 == index ? grid_247 : _GEN_573; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_575 = 9'hf8 == index ? grid_248 : _GEN_574; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_576 = 9'hf9 == index ? grid_249 : _GEN_575; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_577 = 9'hfa == index ? grid_250 : _GEN_576; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_578 = 9'hfb == index ? grid_251 : _GEN_577; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_579 = 9'hfc == index ? grid_252 : _GEN_578; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_580 = 9'hfd == index ? grid_253 : _GEN_579; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_581 = 9'hfe == index ? grid_254 : _GEN_580; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_582 = 9'hff == index ? grid_255 : _GEN_581; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_583 = 9'h100 == index ? grid_256 : _GEN_582; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_584 = 9'h101 == index ? grid_257 : _GEN_583; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_585 = 9'h102 == index ? grid_258 : _GEN_584; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_586 = 9'h103 == index ? grid_259 : _GEN_585; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_587 = 9'h104 == index ? grid_260 : _GEN_586; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_588 = 9'h105 == index ? grid_261 : _GEN_587; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_589 = 9'h106 == index ? grid_262 : _GEN_588; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_590 = 9'h107 == index ? grid_263 : _GEN_589; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_591 = 9'h108 == index ? grid_264 : _GEN_590; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_592 = 9'h109 == index ? grid_265 : _GEN_591; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_593 = 9'h10a == index ? grid_266 : _GEN_592; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_594 = 9'h10b == index ? grid_267 : _GEN_593; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_595 = 9'h10c == index ? grid_268 : _GEN_594; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_596 = 9'h10d == index ? grid_269 : _GEN_595; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_597 = 9'h10e == index ? grid_270 : _GEN_596; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_598 = 9'h10f == index ? grid_271 : _GEN_597; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_599 = 9'h110 == index ? grid_272 : _GEN_598; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_600 = 9'h111 == index ? grid_273 : _GEN_599; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_601 = 9'h112 == index ? grid_274 : _GEN_600; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_602 = 9'h113 == index ? grid_275 : _GEN_601; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_603 = 9'h114 == index ? grid_276 : _GEN_602; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_604 = 9'h115 == index ? grid_277 : _GEN_603; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_605 = 9'h116 == index ? grid_278 : _GEN_604; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_606 = 9'h117 == index ? grid_279 : _GEN_605; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_607 = 9'h118 == index ? grid_280 : _GEN_606; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_608 = 9'h119 == index ? grid_281 : _GEN_607; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_609 = 9'h11a == index ? grid_282 : _GEN_608; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_610 = 9'h11b == index ? grid_283 : _GEN_609; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_611 = 9'h11c == index ? grid_284 : _GEN_610; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_612 = 9'h11d == index ? grid_285 : _GEN_611; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_613 = 9'h11e == index ? grid_286 : _GEN_612; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_614 = 9'h11f == index ? grid_287 : _GEN_613; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_615 = 9'h120 == index ? grid_288 : _GEN_614; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_616 = 9'h121 == index ? grid_289 : _GEN_615; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_617 = 9'h122 == index ? grid_290 : _GEN_616; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_618 = 9'h123 == index ? grid_291 : _GEN_617; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_619 = 9'h124 == index ? grid_292 : _GEN_618; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_620 = 9'h125 == index ? grid_293 : _GEN_619; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_621 = 9'h126 == index ? grid_294 : _GEN_620; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_622 = 9'h127 == index ? grid_295 : _GEN_621; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_623 = 9'h128 == index ? grid_296 : _GEN_622; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_624 = 9'h129 == index ? grid_297 : _GEN_623; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_625 = 9'h12a == index ? grid_298 : _GEN_624; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_626 = 9'h12b == index ? grid_299 : _GEN_625; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_628 = 9'h1 == _aboveValue_T_1 ? grid_1 : grid_0; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_629 = 9'h2 == _aboveValue_T_1 ? grid_2 : _GEN_628; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_630 = 9'h3 == _aboveValue_T_1 ? grid_3 : _GEN_629; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_631 = 9'h4 == _aboveValue_T_1 ? grid_4 : _GEN_630; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_632 = 9'h5 == _aboveValue_T_1 ? grid_5 : _GEN_631; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_633 = 9'h6 == _aboveValue_T_1 ? grid_6 : _GEN_632; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_634 = 9'h7 == _aboveValue_T_1 ? grid_7 : _GEN_633; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_635 = 9'h8 == _aboveValue_T_1 ? grid_8 : _GEN_634; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_636 = 9'h9 == _aboveValue_T_1 ? grid_9 : _GEN_635; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_637 = 9'ha == _aboveValue_T_1 ? grid_10 : _GEN_636; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_638 = 9'hb == _aboveValue_T_1 ? grid_11 : _GEN_637; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_639 = 9'hc == _aboveValue_T_1 ? grid_12 : _GEN_638; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_640 = 9'hd == _aboveValue_T_1 ? grid_13 : _GEN_639; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_641 = 9'he == _aboveValue_T_1 ? grid_14 : _GEN_640; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_642 = 9'hf == _aboveValue_T_1 ? grid_15 : _GEN_641; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_643 = 9'h10 == _aboveValue_T_1 ? grid_16 : _GEN_642; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_644 = 9'h11 == _aboveValue_T_1 ? grid_17 : _GEN_643; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_645 = 9'h12 == _aboveValue_T_1 ? grid_18 : _GEN_644; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_646 = 9'h13 == _aboveValue_T_1 ? grid_19 : _GEN_645; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_647 = 9'h14 == _aboveValue_T_1 ? grid_20 : _GEN_646; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_648 = 9'h15 == _aboveValue_T_1 ? grid_21 : _GEN_647; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_649 = 9'h16 == _aboveValue_T_1 ? grid_22 : _GEN_648; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_650 = 9'h17 == _aboveValue_T_1 ? grid_23 : _GEN_649; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_651 = 9'h18 == _aboveValue_T_1 ? grid_24 : _GEN_650; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_652 = 9'h19 == _aboveValue_T_1 ? grid_25 : _GEN_651; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_653 = 9'h1a == _aboveValue_T_1 ? grid_26 : _GEN_652; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_654 = 9'h1b == _aboveValue_T_1 ? grid_27 : _GEN_653; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_655 = 9'h1c == _aboveValue_T_1 ? grid_28 : _GEN_654; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_656 = 9'h1d == _aboveValue_T_1 ? grid_29 : _GEN_655; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_657 = 9'h1e == _aboveValue_T_1 ? grid_30 : _GEN_656; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_658 = 9'h1f == _aboveValue_T_1 ? grid_31 : _GEN_657; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_659 = 9'h20 == _aboveValue_T_1 ? grid_32 : _GEN_658; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_660 = 9'h21 == _aboveValue_T_1 ? grid_33 : _GEN_659; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_661 = 9'h22 == _aboveValue_T_1 ? grid_34 : _GEN_660; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_662 = 9'h23 == _aboveValue_T_1 ? grid_35 : _GEN_661; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_663 = 9'h24 == _aboveValue_T_1 ? grid_36 : _GEN_662; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_664 = 9'h25 == _aboveValue_T_1 ? grid_37 : _GEN_663; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_665 = 9'h26 == _aboveValue_T_1 ? grid_38 : _GEN_664; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_666 = 9'h27 == _aboveValue_T_1 ? grid_39 : _GEN_665; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_667 = 9'h28 == _aboveValue_T_1 ? grid_40 : _GEN_666; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_668 = 9'h29 == _aboveValue_T_1 ? grid_41 : _GEN_667; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_669 = 9'h2a == _aboveValue_T_1 ? grid_42 : _GEN_668; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_670 = 9'h2b == _aboveValue_T_1 ? grid_43 : _GEN_669; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_671 = 9'h2c == _aboveValue_T_1 ? grid_44 : _GEN_670; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_672 = 9'h2d == _aboveValue_T_1 ? grid_45 : _GEN_671; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_673 = 9'h2e == _aboveValue_T_1 ? grid_46 : _GEN_672; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_674 = 9'h2f == _aboveValue_T_1 ? grid_47 : _GEN_673; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_675 = 9'h30 == _aboveValue_T_1 ? grid_48 : _GEN_674; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_676 = 9'h31 == _aboveValue_T_1 ? grid_49 : _GEN_675; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_677 = 9'h32 == _aboveValue_T_1 ? grid_50 : _GEN_676; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_678 = 9'h33 == _aboveValue_T_1 ? grid_51 : _GEN_677; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_679 = 9'h34 == _aboveValue_T_1 ? grid_52 : _GEN_678; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_680 = 9'h35 == _aboveValue_T_1 ? grid_53 : _GEN_679; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_681 = 9'h36 == _aboveValue_T_1 ? grid_54 : _GEN_680; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_682 = 9'h37 == _aboveValue_T_1 ? grid_55 : _GEN_681; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_683 = 9'h38 == _aboveValue_T_1 ? grid_56 : _GEN_682; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_684 = 9'h39 == _aboveValue_T_1 ? grid_57 : _GEN_683; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_685 = 9'h3a == _aboveValue_T_1 ? grid_58 : _GEN_684; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_686 = 9'h3b == _aboveValue_T_1 ? grid_59 : _GEN_685; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_687 = 9'h3c == _aboveValue_T_1 ? grid_60 : _GEN_686; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_688 = 9'h3d == _aboveValue_T_1 ? grid_61 : _GEN_687; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_689 = 9'h3e == _aboveValue_T_1 ? grid_62 : _GEN_688; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_690 = 9'h3f == _aboveValue_T_1 ? grid_63 : _GEN_689; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_691 = 9'h40 == _aboveValue_T_1 ? grid_64 : _GEN_690; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_692 = 9'h41 == _aboveValue_T_1 ? grid_65 : _GEN_691; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_693 = 9'h42 == _aboveValue_T_1 ? grid_66 : _GEN_692; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_694 = 9'h43 == _aboveValue_T_1 ? grid_67 : _GEN_693; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_695 = 9'h44 == _aboveValue_T_1 ? grid_68 : _GEN_694; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_696 = 9'h45 == _aboveValue_T_1 ? grid_69 : _GEN_695; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_697 = 9'h46 == _aboveValue_T_1 ? grid_70 : _GEN_696; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_698 = 9'h47 == _aboveValue_T_1 ? grid_71 : _GEN_697; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_699 = 9'h48 == _aboveValue_T_1 ? grid_72 : _GEN_698; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_700 = 9'h49 == _aboveValue_T_1 ? grid_73 : _GEN_699; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_701 = 9'h4a == _aboveValue_T_1 ? grid_74 : _GEN_700; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_702 = 9'h4b == _aboveValue_T_1 ? grid_75 : _GEN_701; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_703 = 9'h4c == _aboveValue_T_1 ? grid_76 : _GEN_702; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_704 = 9'h4d == _aboveValue_T_1 ? grid_77 : _GEN_703; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_705 = 9'h4e == _aboveValue_T_1 ? grid_78 : _GEN_704; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_706 = 9'h4f == _aboveValue_T_1 ? grid_79 : _GEN_705; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_707 = 9'h50 == _aboveValue_T_1 ? grid_80 : _GEN_706; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_708 = 9'h51 == _aboveValue_T_1 ? grid_81 : _GEN_707; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_709 = 9'h52 == _aboveValue_T_1 ? grid_82 : _GEN_708; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_710 = 9'h53 == _aboveValue_T_1 ? grid_83 : _GEN_709; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_711 = 9'h54 == _aboveValue_T_1 ? grid_84 : _GEN_710; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_712 = 9'h55 == _aboveValue_T_1 ? grid_85 : _GEN_711; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_713 = 9'h56 == _aboveValue_T_1 ? grid_86 : _GEN_712; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_714 = 9'h57 == _aboveValue_T_1 ? grid_87 : _GEN_713; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_715 = 9'h58 == _aboveValue_T_1 ? grid_88 : _GEN_714; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_716 = 9'h59 == _aboveValue_T_1 ? grid_89 : _GEN_715; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_717 = 9'h5a == _aboveValue_T_1 ? grid_90 : _GEN_716; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_718 = 9'h5b == _aboveValue_T_1 ? grid_91 : _GEN_717; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_719 = 9'h5c == _aboveValue_T_1 ? grid_92 : _GEN_718; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_720 = 9'h5d == _aboveValue_T_1 ? grid_93 : _GEN_719; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_721 = 9'h5e == _aboveValue_T_1 ? grid_94 : _GEN_720; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_722 = 9'h5f == _aboveValue_T_1 ? grid_95 : _GEN_721; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_723 = 9'h60 == _aboveValue_T_1 ? grid_96 : _GEN_722; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_724 = 9'h61 == _aboveValue_T_1 ? grid_97 : _GEN_723; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_725 = 9'h62 == _aboveValue_T_1 ? grid_98 : _GEN_724; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_726 = 9'h63 == _aboveValue_T_1 ? grid_99 : _GEN_725; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_727 = 9'h64 == _aboveValue_T_1 ? grid_100 : _GEN_726; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_728 = 9'h65 == _aboveValue_T_1 ? grid_101 : _GEN_727; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_729 = 9'h66 == _aboveValue_T_1 ? grid_102 : _GEN_728; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_730 = 9'h67 == _aboveValue_T_1 ? grid_103 : _GEN_729; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_731 = 9'h68 == _aboveValue_T_1 ? grid_104 : _GEN_730; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_732 = 9'h69 == _aboveValue_T_1 ? grid_105 : _GEN_731; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_733 = 9'h6a == _aboveValue_T_1 ? grid_106 : _GEN_732; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_734 = 9'h6b == _aboveValue_T_1 ? grid_107 : _GEN_733; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_735 = 9'h6c == _aboveValue_T_1 ? grid_108 : _GEN_734; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_736 = 9'h6d == _aboveValue_T_1 ? grid_109 : _GEN_735; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_737 = 9'h6e == _aboveValue_T_1 ? grid_110 : _GEN_736; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_738 = 9'h6f == _aboveValue_T_1 ? grid_111 : _GEN_737; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_739 = 9'h70 == _aboveValue_T_1 ? grid_112 : _GEN_738; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_740 = 9'h71 == _aboveValue_T_1 ? grid_113 : _GEN_739; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_741 = 9'h72 == _aboveValue_T_1 ? grid_114 : _GEN_740; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_742 = 9'h73 == _aboveValue_T_1 ? grid_115 : _GEN_741; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_743 = 9'h74 == _aboveValue_T_1 ? grid_116 : _GEN_742; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_744 = 9'h75 == _aboveValue_T_1 ? grid_117 : _GEN_743; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_745 = 9'h76 == _aboveValue_T_1 ? grid_118 : _GEN_744; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_746 = 9'h77 == _aboveValue_T_1 ? grid_119 : _GEN_745; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_747 = 9'h78 == _aboveValue_T_1 ? grid_120 : _GEN_746; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_748 = 9'h79 == _aboveValue_T_1 ? grid_121 : _GEN_747; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_749 = 9'h7a == _aboveValue_T_1 ? grid_122 : _GEN_748; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_750 = 9'h7b == _aboveValue_T_1 ? grid_123 : _GEN_749; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_751 = 9'h7c == _aboveValue_T_1 ? grid_124 : _GEN_750; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_752 = 9'h7d == _aboveValue_T_1 ? grid_125 : _GEN_751; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_753 = 9'h7e == _aboveValue_T_1 ? grid_126 : _GEN_752; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_754 = 9'h7f == _aboveValue_T_1 ? grid_127 : _GEN_753; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_755 = 9'h80 == _aboveValue_T_1 ? grid_128 : _GEN_754; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_756 = 9'h81 == _aboveValue_T_1 ? grid_129 : _GEN_755; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_757 = 9'h82 == _aboveValue_T_1 ? grid_130 : _GEN_756; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_758 = 9'h83 == _aboveValue_T_1 ? grid_131 : _GEN_757; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_759 = 9'h84 == _aboveValue_T_1 ? grid_132 : _GEN_758; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_760 = 9'h85 == _aboveValue_T_1 ? grid_133 : _GEN_759; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_761 = 9'h86 == _aboveValue_T_1 ? grid_134 : _GEN_760; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_762 = 9'h87 == _aboveValue_T_1 ? grid_135 : _GEN_761; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_763 = 9'h88 == _aboveValue_T_1 ? grid_136 : _GEN_762; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_764 = 9'h89 == _aboveValue_T_1 ? grid_137 : _GEN_763; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_765 = 9'h8a == _aboveValue_T_1 ? grid_138 : _GEN_764; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_766 = 9'h8b == _aboveValue_T_1 ? grid_139 : _GEN_765; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_767 = 9'h8c == _aboveValue_T_1 ? grid_140 : _GEN_766; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_768 = 9'h8d == _aboveValue_T_1 ? grid_141 : _GEN_767; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_769 = 9'h8e == _aboveValue_T_1 ? grid_142 : _GEN_768; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_770 = 9'h8f == _aboveValue_T_1 ? grid_143 : _GEN_769; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_771 = 9'h90 == _aboveValue_T_1 ? grid_144 : _GEN_770; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_772 = 9'h91 == _aboveValue_T_1 ? grid_145 : _GEN_771; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_773 = 9'h92 == _aboveValue_T_1 ? grid_146 : _GEN_772; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_774 = 9'h93 == _aboveValue_T_1 ? grid_147 : _GEN_773; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_775 = 9'h94 == _aboveValue_T_1 ? grid_148 : _GEN_774; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_776 = 9'h95 == _aboveValue_T_1 ? grid_149 : _GEN_775; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_777 = 9'h96 == _aboveValue_T_1 ? grid_150 : _GEN_776; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_778 = 9'h97 == _aboveValue_T_1 ? grid_151 : _GEN_777; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_779 = 9'h98 == _aboveValue_T_1 ? grid_152 : _GEN_778; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_780 = 9'h99 == _aboveValue_T_1 ? grid_153 : _GEN_779; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_781 = 9'h9a == _aboveValue_T_1 ? grid_154 : _GEN_780; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_782 = 9'h9b == _aboveValue_T_1 ? grid_155 : _GEN_781; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_783 = 9'h9c == _aboveValue_T_1 ? grid_156 : _GEN_782; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_784 = 9'h9d == _aboveValue_T_1 ? grid_157 : _GEN_783; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_785 = 9'h9e == _aboveValue_T_1 ? grid_158 : _GEN_784; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_786 = 9'h9f == _aboveValue_T_1 ? grid_159 : _GEN_785; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_787 = 9'ha0 == _aboveValue_T_1 ? grid_160 : _GEN_786; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_788 = 9'ha1 == _aboveValue_T_1 ? grid_161 : _GEN_787; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_789 = 9'ha2 == _aboveValue_T_1 ? grid_162 : _GEN_788; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_790 = 9'ha3 == _aboveValue_T_1 ? grid_163 : _GEN_789; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_791 = 9'ha4 == _aboveValue_T_1 ? grid_164 : _GEN_790; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_792 = 9'ha5 == _aboveValue_T_1 ? grid_165 : _GEN_791; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_793 = 9'ha6 == _aboveValue_T_1 ? grid_166 : _GEN_792; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_794 = 9'ha7 == _aboveValue_T_1 ? grid_167 : _GEN_793; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_795 = 9'ha8 == _aboveValue_T_1 ? grid_168 : _GEN_794; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_796 = 9'ha9 == _aboveValue_T_1 ? grid_169 : _GEN_795; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_797 = 9'haa == _aboveValue_T_1 ? grid_170 : _GEN_796; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_798 = 9'hab == _aboveValue_T_1 ? grid_171 : _GEN_797; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_799 = 9'hac == _aboveValue_T_1 ? grid_172 : _GEN_798; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_800 = 9'had == _aboveValue_T_1 ? grid_173 : _GEN_799; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_801 = 9'hae == _aboveValue_T_1 ? grid_174 : _GEN_800; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_802 = 9'haf == _aboveValue_T_1 ? grid_175 : _GEN_801; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_803 = 9'hb0 == _aboveValue_T_1 ? grid_176 : _GEN_802; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_804 = 9'hb1 == _aboveValue_T_1 ? grid_177 : _GEN_803; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_805 = 9'hb2 == _aboveValue_T_1 ? grid_178 : _GEN_804; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_806 = 9'hb3 == _aboveValue_T_1 ? grid_179 : _GEN_805; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_807 = 9'hb4 == _aboveValue_T_1 ? grid_180 : _GEN_806; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_808 = 9'hb5 == _aboveValue_T_1 ? grid_181 : _GEN_807; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_809 = 9'hb6 == _aboveValue_T_1 ? grid_182 : _GEN_808; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_810 = 9'hb7 == _aboveValue_T_1 ? grid_183 : _GEN_809; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_811 = 9'hb8 == _aboveValue_T_1 ? grid_184 : _GEN_810; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_812 = 9'hb9 == _aboveValue_T_1 ? grid_185 : _GEN_811; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_813 = 9'hba == _aboveValue_T_1 ? grid_186 : _GEN_812; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_814 = 9'hbb == _aboveValue_T_1 ? grid_187 : _GEN_813; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_815 = 9'hbc == _aboveValue_T_1 ? grid_188 : _GEN_814; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_816 = 9'hbd == _aboveValue_T_1 ? grid_189 : _GEN_815; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_817 = 9'hbe == _aboveValue_T_1 ? grid_190 : _GEN_816; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_818 = 9'hbf == _aboveValue_T_1 ? grid_191 : _GEN_817; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_819 = 9'hc0 == _aboveValue_T_1 ? grid_192 : _GEN_818; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_820 = 9'hc1 == _aboveValue_T_1 ? grid_193 : _GEN_819; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_821 = 9'hc2 == _aboveValue_T_1 ? grid_194 : _GEN_820; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_822 = 9'hc3 == _aboveValue_T_1 ? grid_195 : _GEN_821; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_823 = 9'hc4 == _aboveValue_T_1 ? grid_196 : _GEN_822; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_824 = 9'hc5 == _aboveValue_T_1 ? grid_197 : _GEN_823; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_825 = 9'hc6 == _aboveValue_T_1 ? grid_198 : _GEN_824; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_826 = 9'hc7 == _aboveValue_T_1 ? grid_199 : _GEN_825; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_827 = 9'hc8 == _aboveValue_T_1 ? grid_200 : _GEN_826; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_828 = 9'hc9 == _aboveValue_T_1 ? grid_201 : _GEN_827; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_829 = 9'hca == _aboveValue_T_1 ? grid_202 : _GEN_828; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_830 = 9'hcb == _aboveValue_T_1 ? grid_203 : _GEN_829; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_831 = 9'hcc == _aboveValue_T_1 ? grid_204 : _GEN_830; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_832 = 9'hcd == _aboveValue_T_1 ? grid_205 : _GEN_831; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_833 = 9'hce == _aboveValue_T_1 ? grid_206 : _GEN_832; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_834 = 9'hcf == _aboveValue_T_1 ? grid_207 : _GEN_833; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_835 = 9'hd0 == _aboveValue_T_1 ? grid_208 : _GEN_834; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_836 = 9'hd1 == _aboveValue_T_1 ? grid_209 : _GEN_835; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_837 = 9'hd2 == _aboveValue_T_1 ? grid_210 : _GEN_836; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_838 = 9'hd3 == _aboveValue_T_1 ? grid_211 : _GEN_837; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_839 = 9'hd4 == _aboveValue_T_1 ? grid_212 : _GEN_838; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_840 = 9'hd5 == _aboveValue_T_1 ? grid_213 : _GEN_839; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_841 = 9'hd6 == _aboveValue_T_1 ? grid_214 : _GEN_840; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_842 = 9'hd7 == _aboveValue_T_1 ? grid_215 : _GEN_841; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_843 = 9'hd8 == _aboveValue_T_1 ? grid_216 : _GEN_842; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_844 = 9'hd9 == _aboveValue_T_1 ? grid_217 : _GEN_843; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_845 = 9'hda == _aboveValue_T_1 ? grid_218 : _GEN_844; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_846 = 9'hdb == _aboveValue_T_1 ? grid_219 : _GEN_845; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_847 = 9'hdc == _aboveValue_T_1 ? grid_220 : _GEN_846; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_848 = 9'hdd == _aboveValue_T_1 ? grid_221 : _GEN_847; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_849 = 9'hde == _aboveValue_T_1 ? grid_222 : _GEN_848; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_850 = 9'hdf == _aboveValue_T_1 ? grid_223 : _GEN_849; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_851 = 9'he0 == _aboveValue_T_1 ? grid_224 : _GEN_850; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_852 = 9'he1 == _aboveValue_T_1 ? grid_225 : _GEN_851; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_853 = 9'he2 == _aboveValue_T_1 ? grid_226 : _GEN_852; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_854 = 9'he3 == _aboveValue_T_1 ? grid_227 : _GEN_853; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_855 = 9'he4 == _aboveValue_T_1 ? grid_228 : _GEN_854; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_856 = 9'he5 == _aboveValue_T_1 ? grid_229 : _GEN_855; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_857 = 9'he6 == _aboveValue_T_1 ? grid_230 : _GEN_856; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_858 = 9'he7 == _aboveValue_T_1 ? grid_231 : _GEN_857; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_859 = 9'he8 == _aboveValue_T_1 ? grid_232 : _GEN_858; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_860 = 9'he9 == _aboveValue_T_1 ? grid_233 : _GEN_859; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_861 = 9'hea == _aboveValue_T_1 ? grid_234 : _GEN_860; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_862 = 9'heb == _aboveValue_T_1 ? grid_235 : _GEN_861; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_863 = 9'hec == _aboveValue_T_1 ? grid_236 : _GEN_862; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_864 = 9'hed == _aboveValue_T_1 ? grid_237 : _GEN_863; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_865 = 9'hee == _aboveValue_T_1 ? grid_238 : _GEN_864; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_866 = 9'hef == _aboveValue_T_1 ? grid_239 : _GEN_865; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_867 = 9'hf0 == _aboveValue_T_1 ? grid_240 : _GEN_866; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_868 = 9'hf1 == _aboveValue_T_1 ? grid_241 : _GEN_867; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_869 = 9'hf2 == _aboveValue_T_1 ? grid_242 : _GEN_868; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_870 = 9'hf3 == _aboveValue_T_1 ? grid_243 : _GEN_869; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_871 = 9'hf4 == _aboveValue_T_1 ? grid_244 : _GEN_870; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_872 = 9'hf5 == _aboveValue_T_1 ? grid_245 : _GEN_871; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_873 = 9'hf6 == _aboveValue_T_1 ? grid_246 : _GEN_872; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_874 = 9'hf7 == _aboveValue_T_1 ? grid_247 : _GEN_873; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_875 = 9'hf8 == _aboveValue_T_1 ? grid_248 : _GEN_874; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_876 = 9'hf9 == _aboveValue_T_1 ? grid_249 : _GEN_875; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_877 = 9'hfa == _aboveValue_T_1 ? grid_250 : _GEN_876; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_878 = 9'hfb == _aboveValue_T_1 ? grid_251 : _GEN_877; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_879 = 9'hfc == _aboveValue_T_1 ? grid_252 : _GEN_878; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_880 = 9'hfd == _aboveValue_T_1 ? grid_253 : _GEN_879; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_881 = 9'hfe == _aboveValue_T_1 ? grid_254 : _GEN_880; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_882 = 9'hff == _aboveValue_T_1 ? grid_255 : _GEN_881; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_883 = 9'h100 == _aboveValue_T_1 ? grid_256 : _GEN_882; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_884 = 9'h101 == _aboveValue_T_1 ? grid_257 : _GEN_883; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_885 = 9'h102 == _aboveValue_T_1 ? grid_258 : _GEN_884; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_886 = 9'h103 == _aboveValue_T_1 ? grid_259 : _GEN_885; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_887 = 9'h104 == _aboveValue_T_1 ? grid_260 : _GEN_886; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_888 = 9'h105 == _aboveValue_T_1 ? grid_261 : _GEN_887; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_889 = 9'h106 == _aboveValue_T_1 ? grid_262 : _GEN_888; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_890 = 9'h107 == _aboveValue_T_1 ? grid_263 : _GEN_889; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_891 = 9'h108 == _aboveValue_T_1 ? grid_264 : _GEN_890; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_892 = 9'h109 == _aboveValue_T_1 ? grid_265 : _GEN_891; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_893 = 9'h10a == _aboveValue_T_1 ? grid_266 : _GEN_892; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_894 = 9'h10b == _aboveValue_T_1 ? grid_267 : _GEN_893; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_895 = 9'h10c == _aboveValue_T_1 ? grid_268 : _GEN_894; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_896 = 9'h10d == _aboveValue_T_1 ? grid_269 : _GEN_895; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_897 = 9'h10e == _aboveValue_T_1 ? grid_270 : _GEN_896; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_898 = 9'h10f == _aboveValue_T_1 ? grid_271 : _GEN_897; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_899 = 9'h110 == _aboveValue_T_1 ? grid_272 : _GEN_898; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_900 = 9'h111 == _aboveValue_T_1 ? grid_273 : _GEN_899; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_901 = 9'h112 == _aboveValue_T_1 ? grid_274 : _GEN_900; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_902 = 9'h113 == _aboveValue_T_1 ? grid_275 : _GEN_901; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_903 = 9'h114 == _aboveValue_T_1 ? grid_276 : _GEN_902; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_904 = 9'h115 == _aboveValue_T_1 ? grid_277 : _GEN_903; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_905 = 9'h116 == _aboveValue_T_1 ? grid_278 : _GEN_904; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_906 = 9'h117 == _aboveValue_T_1 ? grid_279 : _GEN_905; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_907 = 9'h118 == _aboveValue_T_1 ? grid_280 : _GEN_906; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_908 = 9'h119 == _aboveValue_T_1 ? grid_281 : _GEN_907; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_909 = 9'h11a == _aboveValue_T_1 ? grid_282 : _GEN_908; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_910 = 9'h11b == _aboveValue_T_1 ? grid_283 : _GEN_909; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_911 = 9'h11c == _aboveValue_T_1 ? grid_284 : _GEN_910; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_912 = 9'h11d == _aboveValue_T_1 ? grid_285 : _GEN_911; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_913 = 9'h11e == _aboveValue_T_1 ? grid_286 : _GEN_912; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_914 = 9'h11f == _aboveValue_T_1 ? grid_287 : _GEN_913; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_915 = 9'h120 == _aboveValue_T_1 ? grid_288 : _GEN_914; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_916 = 9'h121 == _aboveValue_T_1 ? grid_289 : _GEN_915; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_917 = 9'h122 == _aboveValue_T_1 ? grid_290 : _GEN_916; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_918 = 9'h123 == _aboveValue_T_1 ? grid_291 : _GEN_917; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_919 = 9'h124 == _aboveValue_T_1 ? grid_292 : _GEN_918; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_920 = 9'h125 == _aboveValue_T_1 ? grid_293 : _GEN_919; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_921 = 9'h126 == _aboveValue_T_1 ? grid_294 : _GEN_920; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_922 = 9'h127 == _aboveValue_T_1 ? grid_295 : _GEN_921; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_923 = 9'h128 == _aboveValue_T_1 ? grid_296 : _GEN_922; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_924 = 9'h129 == _aboveValue_T_1 ? grid_297 : _GEN_923; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_925 = 9'h12a == _aboveValue_T_1 ? grid_298 : _GEN_924; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [1:0] _GEN_926 = 9'h12b == _aboveValue_T_1 ? grid_299 : _GEN_925; // @[\\src\\main\\scala\\GameLogic.scala 230:{35,35}]
  wire [4:0] _GEN_3496 = {{3'd0}, _GEN_926}; // @[\\src\\main\\scala\\GameLogic.scala 231:46]
  wire [4:0] _io_backBufferWriteData_T_1 = 5'h14 + _GEN_3496; // @[\\src\\main\\scala\\GameLogic.scala 231:46]
  wire [1:0] _GEN_927 = 9'h0 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_928 = 9'h1 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_929 = 9'h2 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_930 = 9'h3 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_931 = 9'h4 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_932 = 9'h5 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_933 = 9'h6 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_934 = 9'h7 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_935 = 9'h8 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_936 = 9'h9 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_937 = 9'ha == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_938 = 9'hb == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_939 = 9'hc == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_940 = 9'hd == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_941 = 9'he == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_942 = 9'hf == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_943 = 9'h10 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_944 = 9'h11 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_945 = 9'h12 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_946 = 9'h13 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_947 = 9'h14 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_948 = 9'h15 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_949 = 9'h16 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_950 = 9'h17 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_951 = 9'h18 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 95:13]
  wire [1:0] _GEN_952 = 9'h19 == index ? _GEN_926 : grid_25; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_953 = 9'h1a == index ? _GEN_926 : grid_26; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_954 = 9'h1b == index ? _GEN_926 : grid_27; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_955 = 9'h1c == index ? _GEN_926 : grid_28; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_956 = 9'h1d == index ? _GEN_926 : grid_29; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_957 = 9'h1e == index ? _GEN_926 : grid_30; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_958 = 9'h1f == index ? _GEN_926 : grid_31; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_959 = 9'h20 == index ? _GEN_926 : grid_32; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_960 = 9'h21 == index ? _GEN_926 : grid_33; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_961 = 9'h22 == index ? _GEN_926 : grid_34; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_962 = 9'h23 == index ? _GEN_926 : grid_35; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_963 = 9'h24 == index ? _GEN_926 : grid_36; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_964 = 9'h25 == index ? _GEN_926 : grid_37; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_965 = 9'h26 == index ? _GEN_926 : grid_38; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_966 = 9'h27 == index ? _GEN_926 : grid_39; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_967 = 9'h28 == index ? _GEN_926 : grid_40; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_968 = 9'h29 == index ? _GEN_926 : grid_41; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_969 = 9'h2a == index ? _GEN_926 : grid_42; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_970 = 9'h2b == index ? _GEN_926 : grid_43; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_971 = 9'h2c == index ? _GEN_926 : grid_44; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_972 = 9'h2d == index ? _GEN_926 : grid_45; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_973 = 9'h2e == index ? _GEN_926 : grid_46; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_974 = 9'h2f == index ? _GEN_926 : grid_47; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_975 = 9'h30 == index ? _GEN_926 : grid_48; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_976 = 9'h31 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_977 = 9'h32 == index ? _GEN_926 : grid_50; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_978 = 9'h33 == index ? _GEN_926 : grid_51; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_979 = 9'h34 == index ? _GEN_926 : grid_52; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_980 = 9'h35 == index ? _GEN_926 : grid_53; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_981 = 9'h36 == index ? _GEN_926 : grid_54; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_982 = 9'h37 == index ? _GEN_926 : grid_55; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_983 = 9'h38 == index ? _GEN_926 : grid_56; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_984 = 9'h39 == index ? _GEN_926 : grid_57; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_985 = 9'h3a == index ? _GEN_926 : grid_58; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_986 = 9'h3b == index ? _GEN_926 : grid_59; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_987 = 9'h3c == index ? _GEN_926 : grid_60; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_988 = 9'h3d == index ? _GEN_926 : grid_61; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_989 = 9'h3e == index ? _GEN_926 : grid_62; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_990 = 9'h3f == index ? _GEN_926 : grid_63; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_991 = 9'h40 == index ? _GEN_926 : grid_64; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_992 = 9'h41 == index ? _GEN_926 : grid_65; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_993 = 9'h42 == index ? _GEN_926 : grid_66; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_994 = 9'h43 == index ? _GEN_926 : grid_67; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_995 = 9'h44 == index ? _GEN_926 : grid_68; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_996 = 9'h45 == index ? _GEN_926 : grid_69; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_997 = 9'h46 == index ? _GEN_926 : grid_70; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_998 = 9'h47 == index ? _GEN_926 : grid_71; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_999 = 9'h48 == index ? _GEN_926 : grid_72; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1000 = 9'h49 == index ? _GEN_926 : grid_73; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1001 = 9'h4a == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_1002 = 9'h4b == index ? _GEN_926 : grid_75; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1003 = 9'h4c == index ? _GEN_926 : grid_76; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1004 = 9'h4d == index ? _GEN_926 : grid_77; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1005 = 9'h4e == index ? _GEN_926 : grid_78; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1006 = 9'h4f == index ? _GEN_926 : grid_79; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1007 = 9'h50 == index ? _GEN_926 : grid_80; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1008 = 9'h51 == index ? _GEN_926 : grid_81; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1009 = 9'h52 == index ? _GEN_926 : grid_82; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1010 = 9'h53 == index ? _GEN_926 : grid_83; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1011 = 9'h54 == index ? _GEN_926 : grid_84; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1012 = 9'h55 == index ? _GEN_926 : grid_85; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1013 = 9'h56 == index ? _GEN_926 : grid_86; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1014 = 9'h57 == index ? _GEN_926 : grid_87; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1015 = 9'h58 == index ? _GEN_926 : grid_88; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1016 = 9'h59 == index ? _GEN_926 : grid_89; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1017 = 9'h5a == index ? _GEN_926 : grid_90; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1018 = 9'h5b == index ? _GEN_926 : grid_91; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1019 = 9'h5c == index ? _GEN_926 : grid_92; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1020 = 9'h5d == index ? _GEN_926 : grid_93; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1021 = 9'h5e == index ? _GEN_926 : grid_94; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1022 = 9'h5f == index ? _GEN_926 : grid_95; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1023 = 9'h60 == index ? _GEN_926 : grid_96; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1024 = 9'h61 == index ? _GEN_926 : grid_97; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1025 = 9'h62 == index ? _GEN_926 : grid_98; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1026 = 9'h63 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_1027 = 9'h64 == index ? _GEN_926 : grid_100; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1028 = 9'h65 == index ? _GEN_926 : grid_101; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1029 = 9'h66 == index ? _GEN_926 : grid_102; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1030 = 9'h67 == index ? _GEN_926 : grid_103; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1031 = 9'h68 == index ? _GEN_926 : grid_104; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1032 = 9'h69 == index ? _GEN_926 : grid_105; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1033 = 9'h6a == index ? _GEN_926 : grid_106; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1034 = 9'h6b == index ? _GEN_926 : grid_107; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1035 = 9'h6c == index ? _GEN_926 : grid_108; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1036 = 9'h6d == index ? _GEN_926 : grid_109; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1037 = 9'h6e == index ? _GEN_926 : grid_110; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1038 = 9'h6f == index ? _GEN_926 : grid_111; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1039 = 9'h70 == index ? _GEN_926 : grid_112; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1040 = 9'h71 == index ? _GEN_926 : grid_113; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1041 = 9'h72 == index ? _GEN_926 : grid_114; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1042 = 9'h73 == index ? _GEN_926 : grid_115; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1043 = 9'h74 == index ? _GEN_926 : grid_116; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1044 = 9'h75 == index ? _GEN_926 : grid_117; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1045 = 9'h76 == index ? _GEN_926 : grid_118; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1046 = 9'h77 == index ? _GEN_926 : grid_119; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1047 = 9'h78 == index ? _GEN_926 : grid_120; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1048 = 9'h79 == index ? _GEN_926 : grid_121; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1049 = 9'h7a == index ? _GEN_926 : grid_122; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1050 = 9'h7b == index ? _GEN_926 : grid_123; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1051 = 9'h7c == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_1052 = 9'h7d == index ? _GEN_926 : grid_125; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1053 = 9'h7e == index ? _GEN_926 : grid_126; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1054 = 9'h7f == index ? _GEN_926 : grid_127; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1055 = 9'h80 == index ? _GEN_926 : grid_128; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1056 = 9'h81 == index ? _GEN_926 : grid_129; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1057 = 9'h82 == index ? _GEN_926 : grid_130; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1058 = 9'h83 == index ? _GEN_926 : grid_131; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1059 = 9'h84 == index ? _GEN_926 : grid_132; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1060 = 9'h85 == index ? _GEN_926 : grid_133; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1061 = 9'h86 == index ? _GEN_926 : grid_134; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1062 = 9'h87 == index ? _GEN_926 : grid_135; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1063 = 9'h88 == index ? _GEN_926 : grid_136; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1064 = 9'h89 == index ? _GEN_926 : grid_137; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1065 = 9'h8a == index ? _GEN_926 : grid_138; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1066 = 9'h8b == index ? _GEN_926 : grid_139; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1067 = 9'h8c == index ? _GEN_926 : grid_140; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1068 = 9'h8d == index ? _GEN_926 : grid_141; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1069 = 9'h8e == index ? _GEN_926 : grid_142; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1070 = 9'h8f == index ? _GEN_926 : grid_143; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1071 = 9'h90 == index ? _GEN_926 : grid_144; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1072 = 9'h91 == index ? _GEN_926 : grid_145; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1073 = 9'h92 == index ? _GEN_926 : grid_146; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1074 = 9'h93 == index ? _GEN_926 : grid_147; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1075 = 9'h94 == index ? _GEN_926 : grid_148; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1076 = 9'h95 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_1077 = 9'h96 == index ? _GEN_926 : grid_150; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1078 = 9'h97 == index ? _GEN_926 : grid_151; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1079 = 9'h98 == index ? _GEN_926 : grid_152; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1080 = 9'h99 == index ? _GEN_926 : grid_153; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1081 = 9'h9a == index ? _GEN_926 : grid_154; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1082 = 9'h9b == index ? _GEN_926 : grid_155; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1083 = 9'h9c == index ? _GEN_926 : grid_156; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1084 = 9'h9d == index ? _GEN_926 : grid_157; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1085 = 9'h9e == index ? _GEN_926 : grid_158; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1086 = 9'h9f == index ? _GEN_926 : grid_159; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1087 = 9'ha0 == index ? _GEN_926 : grid_160; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1088 = 9'ha1 == index ? _GEN_926 : grid_161; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1089 = 9'ha2 == index ? _GEN_926 : grid_162; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1090 = 9'ha3 == index ? _GEN_926 : grid_163; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1091 = 9'ha4 == index ? _GEN_926 : grid_164; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1092 = 9'ha5 == index ? _GEN_926 : grid_165; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1093 = 9'ha6 == index ? _GEN_926 : grid_166; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1094 = 9'ha7 == index ? _GEN_926 : grid_167; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1095 = 9'ha8 == index ? _GEN_926 : grid_168; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1096 = 9'ha9 == index ? _GEN_926 : grid_169; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1097 = 9'haa == index ? _GEN_926 : grid_170; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1098 = 9'hab == index ? _GEN_926 : grid_171; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1099 = 9'hac == index ? _GEN_926 : grid_172; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1100 = 9'had == index ? _GEN_926 : grid_173; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1101 = 9'hae == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_1102 = 9'haf == index ? _GEN_926 : grid_175; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1103 = 9'hb0 == index ? _GEN_926 : grid_176; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1104 = 9'hb1 == index ? _GEN_926 : grid_177; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1105 = 9'hb2 == index ? _GEN_926 : grid_178; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1106 = 9'hb3 == index ? _GEN_926 : grid_179; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1107 = 9'hb4 == index ? _GEN_926 : grid_180; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1108 = 9'hb5 == index ? _GEN_926 : grid_181; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1109 = 9'hb6 == index ? _GEN_926 : grid_182; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1110 = 9'hb7 == index ? _GEN_926 : grid_183; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1111 = 9'hb8 == index ? _GEN_926 : grid_184; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1112 = 9'hb9 == index ? _GEN_926 : grid_185; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1113 = 9'hba == index ? _GEN_926 : grid_186; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1114 = 9'hbb == index ? _GEN_926 : grid_187; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1115 = 9'hbc == index ? _GEN_926 : grid_188; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1116 = 9'hbd == index ? _GEN_926 : grid_189; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1117 = 9'hbe == index ? _GEN_926 : grid_190; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1118 = 9'hbf == index ? _GEN_926 : grid_191; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1119 = 9'hc0 == index ? _GEN_926 : grid_192; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1120 = 9'hc1 == index ? _GEN_926 : grid_193; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1121 = 9'hc2 == index ? _GEN_926 : grid_194; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1122 = 9'hc3 == index ? _GEN_926 : grid_195; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1123 = 9'hc4 == index ? _GEN_926 : grid_196; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1124 = 9'hc5 == index ? _GEN_926 : grid_197; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1125 = 9'hc6 == index ? _GEN_926 : grid_198; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1126 = 9'hc7 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_1127 = 9'hc8 == index ? _GEN_926 : grid_200; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1128 = 9'hc9 == index ? _GEN_926 : grid_201; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1129 = 9'hca == index ? _GEN_926 : grid_202; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1130 = 9'hcb == index ? _GEN_926 : grid_203; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1131 = 9'hcc == index ? _GEN_926 : grid_204; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1132 = 9'hcd == index ? _GEN_926 : grid_205; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1133 = 9'hce == index ? _GEN_926 : grid_206; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1134 = 9'hcf == index ? _GEN_926 : grid_207; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1135 = 9'hd0 == index ? _GEN_926 : grid_208; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1136 = 9'hd1 == index ? _GEN_926 : grid_209; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1137 = 9'hd2 == index ? _GEN_926 : grid_210; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1138 = 9'hd3 == index ? _GEN_926 : grid_211; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1139 = 9'hd4 == index ? _GEN_926 : grid_212; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1140 = 9'hd5 == index ? _GEN_926 : grid_213; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1141 = 9'hd6 == index ? _GEN_926 : grid_214; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1142 = 9'hd7 == index ? _GEN_926 : grid_215; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1143 = 9'hd8 == index ? _GEN_926 : grid_216; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1144 = 9'hd9 == index ? _GEN_926 : grid_217; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1145 = 9'hda == index ? _GEN_926 : grid_218; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1146 = 9'hdb == index ? _GEN_926 : grid_219; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1147 = 9'hdc == index ? _GEN_926 : grid_220; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1148 = 9'hdd == index ? _GEN_926 : grid_221; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1149 = 9'hde == index ? _GEN_926 : grid_222; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1150 = 9'hdf == index ? _GEN_926 : grid_223; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1151 = 9'he0 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_1152 = 9'he1 == index ? _GEN_926 : grid_225; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1153 = 9'he2 == index ? _GEN_926 : grid_226; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1154 = 9'he3 == index ? _GEN_926 : grid_227; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1155 = 9'he4 == index ? _GEN_926 : grid_228; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1156 = 9'he5 == index ? _GEN_926 : grid_229; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1157 = 9'he6 == index ? _GEN_926 : grid_230; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1158 = 9'he7 == index ? _GEN_926 : grid_231; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1159 = 9'he8 == index ? _GEN_926 : grid_232; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1160 = 9'he9 == index ? _GEN_926 : grid_233; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1161 = 9'hea == index ? _GEN_926 : grid_234; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1162 = 9'heb == index ? _GEN_926 : grid_235; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1163 = 9'hec == index ? _GEN_926 : grid_236; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1164 = 9'hed == index ? _GEN_926 : grid_237; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1165 = 9'hee == index ? _GEN_926 : grid_238; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1166 = 9'hef == index ? _GEN_926 : grid_239; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1167 = 9'hf0 == index ? _GEN_926 : grid_240; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1168 = 9'hf1 == index ? _GEN_926 : grid_241; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1169 = 9'hf2 == index ? _GEN_926 : grid_242; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1170 = 9'hf3 == index ? _GEN_926 : grid_243; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1171 = 9'hf4 == index ? _GEN_926 : grid_244; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1172 = 9'hf5 == index ? _GEN_926 : grid_245; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1173 = 9'hf6 == index ? _GEN_926 : grid_246; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1174 = 9'hf7 == index ? _GEN_926 : grid_247; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1175 = 9'hf8 == index ? _GEN_926 : grid_248; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1176 = 9'hf9 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_1177 = 9'hfa == index ? _GEN_926 : grid_250; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1178 = 9'hfb == index ? _GEN_926 : grid_251; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1179 = 9'hfc == index ? _GEN_926 : grid_252; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1180 = 9'hfd == index ? _GEN_926 : grid_253; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1181 = 9'hfe == index ? _GEN_926 : grid_254; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1182 = 9'hff == index ? _GEN_926 : grid_255; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1183 = 9'h100 == index ? _GEN_926 : grid_256; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1184 = 9'h101 == index ? _GEN_926 : grid_257; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1185 = 9'h102 == index ? _GEN_926 : grid_258; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1186 = 9'h103 == index ? _GEN_926 : grid_259; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1187 = 9'h104 == index ? _GEN_926 : grid_260; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1188 = 9'h105 == index ? _GEN_926 : grid_261; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1189 = 9'h106 == index ? _GEN_926 : grid_262; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1190 = 9'h107 == index ? _GEN_926 : grid_263; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1191 = 9'h108 == index ? _GEN_926 : grid_264; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1192 = 9'h109 == index ? _GEN_926 : grid_265; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1193 = 9'h10a == index ? _GEN_926 : grid_266; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1194 = 9'h10b == index ? _GEN_926 : grid_267; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1195 = 9'h10c == index ? _GEN_926 : grid_268; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1196 = 9'h10d == index ? _GEN_926 : grid_269; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1197 = 9'h10e == index ? _GEN_926 : grid_270; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1198 = 9'h10f == index ? _GEN_926 : grid_271; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1199 = 9'h110 == index ? _GEN_926 : grid_272; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1200 = 9'h111 == index ? _GEN_926 : grid_273; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 88:21]
  wire [1:0] _GEN_1201 = 9'h112 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 91:23]
  wire [1:0] _GEN_1202 = 9'h113 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1203 = 9'h114 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1204 = 9'h115 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1205 = 9'h116 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1206 = 9'h117 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1207 = 9'h118 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1208 = 9'h119 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1209 = 9'h11a == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1210 = 9'h11b == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1211 = 9'h11c == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1212 = 9'h11d == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1213 = 9'h11e == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1214 = 9'h11f == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1215 = 9'h120 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1216 = 9'h121 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1217 = 9'h122 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1218 = 9'h123 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1219 = 9'h124 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1220 = 9'h125 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1221 = 9'h126 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1222 = 9'h127 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1223 = 9'h128 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1224 = 9'h129 == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1225 = 9'h12a == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [1:0] _GEN_1226 = 9'h12b == index ? _GEN_926 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 232:{27,27} 96:21]
  wire [4:0] _GEN_1527 = ~(_GEN_626 == _GEN_926) ? _io_backBufferWriteData_T_1 : 5'h0; // @[\\src\\main\\scala\\GameLogic.scala 128:26 230:53 231:38]
  wire [1:0] _GEN_1528 = ~(_GEN_626 == _GEN_926) ? _GEN_927 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1529 = ~(_GEN_626 == _GEN_926) ? _GEN_928 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1530 = ~(_GEN_626 == _GEN_926) ? _GEN_929 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1531 = ~(_GEN_626 == _GEN_926) ? _GEN_930 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1532 = ~(_GEN_626 == _GEN_926) ? _GEN_931 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1533 = ~(_GEN_626 == _GEN_926) ? _GEN_932 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1534 = ~(_GEN_626 == _GEN_926) ? _GEN_933 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1535 = ~(_GEN_626 == _GEN_926) ? _GEN_934 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1536 = ~(_GEN_626 == _GEN_926) ? _GEN_935 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1537 = ~(_GEN_626 == _GEN_926) ? _GEN_936 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1538 = ~(_GEN_626 == _GEN_926) ? _GEN_937 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1539 = ~(_GEN_626 == _GEN_926) ? _GEN_938 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1540 = ~(_GEN_626 == _GEN_926) ? _GEN_939 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1541 = ~(_GEN_626 == _GEN_926) ? _GEN_940 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1542 = ~(_GEN_626 == _GEN_926) ? _GEN_941 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1543 = ~(_GEN_626 == _GEN_926) ? _GEN_942 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1544 = ~(_GEN_626 == _GEN_926) ? _GEN_943 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1545 = ~(_GEN_626 == _GEN_926) ? _GEN_944 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1546 = ~(_GEN_626 == _GEN_926) ? _GEN_945 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1547 = ~(_GEN_626 == _GEN_926) ? _GEN_946 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1548 = ~(_GEN_626 == _GEN_926) ? _GEN_947 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1549 = ~(_GEN_626 == _GEN_926) ? _GEN_948 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1550 = ~(_GEN_626 == _GEN_926) ? _GEN_949 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1551 = ~(_GEN_626 == _GEN_926) ? _GEN_950 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1552 = ~(_GEN_626 == _GEN_926) ? _GEN_951 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 95:13]
  wire [1:0] _GEN_1553 = ~(_GEN_626 == _GEN_926) ? _GEN_952 : grid_25; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1554 = ~(_GEN_626 == _GEN_926) ? _GEN_953 : grid_26; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1555 = ~(_GEN_626 == _GEN_926) ? _GEN_954 : grid_27; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1556 = ~(_GEN_626 == _GEN_926) ? _GEN_955 : grid_28; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1557 = ~(_GEN_626 == _GEN_926) ? _GEN_956 : grid_29; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1558 = ~(_GEN_626 == _GEN_926) ? _GEN_957 : grid_30; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1559 = ~(_GEN_626 == _GEN_926) ? _GEN_958 : grid_31; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1560 = ~(_GEN_626 == _GEN_926) ? _GEN_959 : grid_32; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1561 = ~(_GEN_626 == _GEN_926) ? _GEN_960 : grid_33; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1562 = ~(_GEN_626 == _GEN_926) ? _GEN_961 : grid_34; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1563 = ~(_GEN_626 == _GEN_926) ? _GEN_962 : grid_35; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1564 = ~(_GEN_626 == _GEN_926) ? _GEN_963 : grid_36; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1565 = ~(_GEN_626 == _GEN_926) ? _GEN_964 : grid_37; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1566 = ~(_GEN_626 == _GEN_926) ? _GEN_965 : grid_38; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1567 = ~(_GEN_626 == _GEN_926) ? _GEN_966 : grid_39; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1568 = ~(_GEN_626 == _GEN_926) ? _GEN_967 : grid_40; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1569 = ~(_GEN_626 == _GEN_926) ? _GEN_968 : grid_41; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1570 = ~(_GEN_626 == _GEN_926) ? _GEN_969 : grid_42; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1571 = ~(_GEN_626 == _GEN_926) ? _GEN_970 : grid_43; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1572 = ~(_GEN_626 == _GEN_926) ? _GEN_971 : grid_44; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1573 = ~(_GEN_626 == _GEN_926) ? _GEN_972 : grid_45; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1574 = ~(_GEN_626 == _GEN_926) ? _GEN_973 : grid_46; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1575 = ~(_GEN_626 == _GEN_926) ? _GEN_974 : grid_47; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1576 = ~(_GEN_626 == _GEN_926) ? _GEN_975 : grid_48; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1577 = ~(_GEN_626 == _GEN_926) ? _GEN_976 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1578 = ~(_GEN_626 == _GEN_926) ? _GEN_977 : grid_50; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1579 = ~(_GEN_626 == _GEN_926) ? _GEN_978 : grid_51; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1580 = ~(_GEN_626 == _GEN_926) ? _GEN_979 : grid_52; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1581 = ~(_GEN_626 == _GEN_926) ? _GEN_980 : grid_53; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1582 = ~(_GEN_626 == _GEN_926) ? _GEN_981 : grid_54; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1583 = ~(_GEN_626 == _GEN_926) ? _GEN_982 : grid_55; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1584 = ~(_GEN_626 == _GEN_926) ? _GEN_983 : grid_56; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1585 = ~(_GEN_626 == _GEN_926) ? _GEN_984 : grid_57; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1586 = ~(_GEN_626 == _GEN_926) ? _GEN_985 : grid_58; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1587 = ~(_GEN_626 == _GEN_926) ? _GEN_986 : grid_59; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1588 = ~(_GEN_626 == _GEN_926) ? _GEN_987 : grid_60; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1589 = ~(_GEN_626 == _GEN_926) ? _GEN_988 : grid_61; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1590 = ~(_GEN_626 == _GEN_926) ? _GEN_989 : grid_62; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1591 = ~(_GEN_626 == _GEN_926) ? _GEN_990 : grid_63; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1592 = ~(_GEN_626 == _GEN_926) ? _GEN_991 : grid_64; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1593 = ~(_GEN_626 == _GEN_926) ? _GEN_992 : grid_65; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1594 = ~(_GEN_626 == _GEN_926) ? _GEN_993 : grid_66; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1595 = ~(_GEN_626 == _GEN_926) ? _GEN_994 : grid_67; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1596 = ~(_GEN_626 == _GEN_926) ? _GEN_995 : grid_68; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1597 = ~(_GEN_626 == _GEN_926) ? _GEN_996 : grid_69; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1598 = ~(_GEN_626 == _GEN_926) ? _GEN_997 : grid_70; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1599 = ~(_GEN_626 == _GEN_926) ? _GEN_998 : grid_71; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1600 = ~(_GEN_626 == _GEN_926) ? _GEN_999 : grid_72; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1601 = ~(_GEN_626 == _GEN_926) ? _GEN_1000 : grid_73; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1602 = ~(_GEN_626 == _GEN_926) ? _GEN_1001 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1603 = ~(_GEN_626 == _GEN_926) ? _GEN_1002 : grid_75; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1604 = ~(_GEN_626 == _GEN_926) ? _GEN_1003 : grid_76; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1605 = ~(_GEN_626 == _GEN_926) ? _GEN_1004 : grid_77; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1606 = ~(_GEN_626 == _GEN_926) ? _GEN_1005 : grid_78; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1607 = ~(_GEN_626 == _GEN_926) ? _GEN_1006 : grid_79; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1608 = ~(_GEN_626 == _GEN_926) ? _GEN_1007 : grid_80; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1609 = ~(_GEN_626 == _GEN_926) ? _GEN_1008 : grid_81; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1610 = ~(_GEN_626 == _GEN_926) ? _GEN_1009 : grid_82; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1611 = ~(_GEN_626 == _GEN_926) ? _GEN_1010 : grid_83; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1612 = ~(_GEN_626 == _GEN_926) ? _GEN_1011 : grid_84; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1613 = ~(_GEN_626 == _GEN_926) ? _GEN_1012 : grid_85; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1614 = ~(_GEN_626 == _GEN_926) ? _GEN_1013 : grid_86; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1615 = ~(_GEN_626 == _GEN_926) ? _GEN_1014 : grid_87; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1616 = ~(_GEN_626 == _GEN_926) ? _GEN_1015 : grid_88; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1617 = ~(_GEN_626 == _GEN_926) ? _GEN_1016 : grid_89; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1618 = ~(_GEN_626 == _GEN_926) ? _GEN_1017 : grid_90; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1619 = ~(_GEN_626 == _GEN_926) ? _GEN_1018 : grid_91; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1620 = ~(_GEN_626 == _GEN_926) ? _GEN_1019 : grid_92; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1621 = ~(_GEN_626 == _GEN_926) ? _GEN_1020 : grid_93; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1622 = ~(_GEN_626 == _GEN_926) ? _GEN_1021 : grid_94; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1623 = ~(_GEN_626 == _GEN_926) ? _GEN_1022 : grid_95; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1624 = ~(_GEN_626 == _GEN_926) ? _GEN_1023 : grid_96; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1625 = ~(_GEN_626 == _GEN_926) ? _GEN_1024 : grid_97; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1626 = ~(_GEN_626 == _GEN_926) ? _GEN_1025 : grid_98; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1627 = ~(_GEN_626 == _GEN_926) ? _GEN_1026 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1628 = ~(_GEN_626 == _GEN_926) ? _GEN_1027 : grid_100; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1629 = ~(_GEN_626 == _GEN_926) ? _GEN_1028 : grid_101; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1630 = ~(_GEN_626 == _GEN_926) ? _GEN_1029 : grid_102; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1631 = ~(_GEN_626 == _GEN_926) ? _GEN_1030 : grid_103; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1632 = ~(_GEN_626 == _GEN_926) ? _GEN_1031 : grid_104; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1633 = ~(_GEN_626 == _GEN_926) ? _GEN_1032 : grid_105; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1634 = ~(_GEN_626 == _GEN_926) ? _GEN_1033 : grid_106; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1635 = ~(_GEN_626 == _GEN_926) ? _GEN_1034 : grid_107; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1636 = ~(_GEN_626 == _GEN_926) ? _GEN_1035 : grid_108; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1637 = ~(_GEN_626 == _GEN_926) ? _GEN_1036 : grid_109; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1638 = ~(_GEN_626 == _GEN_926) ? _GEN_1037 : grid_110; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1639 = ~(_GEN_626 == _GEN_926) ? _GEN_1038 : grid_111; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1640 = ~(_GEN_626 == _GEN_926) ? _GEN_1039 : grid_112; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1641 = ~(_GEN_626 == _GEN_926) ? _GEN_1040 : grid_113; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1642 = ~(_GEN_626 == _GEN_926) ? _GEN_1041 : grid_114; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1643 = ~(_GEN_626 == _GEN_926) ? _GEN_1042 : grid_115; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1644 = ~(_GEN_626 == _GEN_926) ? _GEN_1043 : grid_116; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1645 = ~(_GEN_626 == _GEN_926) ? _GEN_1044 : grid_117; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1646 = ~(_GEN_626 == _GEN_926) ? _GEN_1045 : grid_118; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1647 = ~(_GEN_626 == _GEN_926) ? _GEN_1046 : grid_119; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1648 = ~(_GEN_626 == _GEN_926) ? _GEN_1047 : grid_120; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1649 = ~(_GEN_626 == _GEN_926) ? _GEN_1048 : grid_121; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1650 = ~(_GEN_626 == _GEN_926) ? _GEN_1049 : grid_122; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1651 = ~(_GEN_626 == _GEN_926) ? _GEN_1050 : grid_123; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1652 = ~(_GEN_626 == _GEN_926) ? _GEN_1051 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1653 = ~(_GEN_626 == _GEN_926) ? _GEN_1052 : grid_125; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1654 = ~(_GEN_626 == _GEN_926) ? _GEN_1053 : grid_126; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1655 = ~(_GEN_626 == _GEN_926) ? _GEN_1054 : grid_127; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1656 = ~(_GEN_626 == _GEN_926) ? _GEN_1055 : grid_128; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1657 = ~(_GEN_626 == _GEN_926) ? _GEN_1056 : grid_129; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1658 = ~(_GEN_626 == _GEN_926) ? _GEN_1057 : grid_130; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1659 = ~(_GEN_626 == _GEN_926) ? _GEN_1058 : grid_131; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1660 = ~(_GEN_626 == _GEN_926) ? _GEN_1059 : grid_132; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1661 = ~(_GEN_626 == _GEN_926) ? _GEN_1060 : grid_133; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1662 = ~(_GEN_626 == _GEN_926) ? _GEN_1061 : grid_134; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1663 = ~(_GEN_626 == _GEN_926) ? _GEN_1062 : grid_135; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1664 = ~(_GEN_626 == _GEN_926) ? _GEN_1063 : grid_136; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1665 = ~(_GEN_626 == _GEN_926) ? _GEN_1064 : grid_137; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1666 = ~(_GEN_626 == _GEN_926) ? _GEN_1065 : grid_138; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1667 = ~(_GEN_626 == _GEN_926) ? _GEN_1066 : grid_139; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1668 = ~(_GEN_626 == _GEN_926) ? _GEN_1067 : grid_140; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1669 = ~(_GEN_626 == _GEN_926) ? _GEN_1068 : grid_141; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1670 = ~(_GEN_626 == _GEN_926) ? _GEN_1069 : grid_142; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1671 = ~(_GEN_626 == _GEN_926) ? _GEN_1070 : grid_143; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1672 = ~(_GEN_626 == _GEN_926) ? _GEN_1071 : grid_144; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1673 = ~(_GEN_626 == _GEN_926) ? _GEN_1072 : grid_145; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1674 = ~(_GEN_626 == _GEN_926) ? _GEN_1073 : grid_146; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1675 = ~(_GEN_626 == _GEN_926) ? _GEN_1074 : grid_147; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1676 = ~(_GEN_626 == _GEN_926) ? _GEN_1075 : grid_148; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1677 = ~(_GEN_626 == _GEN_926) ? _GEN_1076 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1678 = ~(_GEN_626 == _GEN_926) ? _GEN_1077 : grid_150; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1679 = ~(_GEN_626 == _GEN_926) ? _GEN_1078 : grid_151; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1680 = ~(_GEN_626 == _GEN_926) ? _GEN_1079 : grid_152; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1681 = ~(_GEN_626 == _GEN_926) ? _GEN_1080 : grid_153; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1682 = ~(_GEN_626 == _GEN_926) ? _GEN_1081 : grid_154; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1683 = ~(_GEN_626 == _GEN_926) ? _GEN_1082 : grid_155; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1684 = ~(_GEN_626 == _GEN_926) ? _GEN_1083 : grid_156; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1685 = ~(_GEN_626 == _GEN_926) ? _GEN_1084 : grid_157; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1686 = ~(_GEN_626 == _GEN_926) ? _GEN_1085 : grid_158; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1687 = ~(_GEN_626 == _GEN_926) ? _GEN_1086 : grid_159; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1688 = ~(_GEN_626 == _GEN_926) ? _GEN_1087 : grid_160; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1689 = ~(_GEN_626 == _GEN_926) ? _GEN_1088 : grid_161; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1690 = ~(_GEN_626 == _GEN_926) ? _GEN_1089 : grid_162; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1691 = ~(_GEN_626 == _GEN_926) ? _GEN_1090 : grid_163; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1692 = ~(_GEN_626 == _GEN_926) ? _GEN_1091 : grid_164; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1693 = ~(_GEN_626 == _GEN_926) ? _GEN_1092 : grid_165; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1694 = ~(_GEN_626 == _GEN_926) ? _GEN_1093 : grid_166; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1695 = ~(_GEN_626 == _GEN_926) ? _GEN_1094 : grid_167; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1696 = ~(_GEN_626 == _GEN_926) ? _GEN_1095 : grid_168; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1697 = ~(_GEN_626 == _GEN_926) ? _GEN_1096 : grid_169; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1698 = ~(_GEN_626 == _GEN_926) ? _GEN_1097 : grid_170; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1699 = ~(_GEN_626 == _GEN_926) ? _GEN_1098 : grid_171; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1700 = ~(_GEN_626 == _GEN_926) ? _GEN_1099 : grid_172; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1701 = ~(_GEN_626 == _GEN_926) ? _GEN_1100 : grid_173; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1702 = ~(_GEN_626 == _GEN_926) ? _GEN_1101 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1703 = ~(_GEN_626 == _GEN_926) ? _GEN_1102 : grid_175; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1704 = ~(_GEN_626 == _GEN_926) ? _GEN_1103 : grid_176; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1705 = ~(_GEN_626 == _GEN_926) ? _GEN_1104 : grid_177; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1706 = ~(_GEN_626 == _GEN_926) ? _GEN_1105 : grid_178; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1707 = ~(_GEN_626 == _GEN_926) ? _GEN_1106 : grid_179; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1708 = ~(_GEN_626 == _GEN_926) ? _GEN_1107 : grid_180; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1709 = ~(_GEN_626 == _GEN_926) ? _GEN_1108 : grid_181; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1710 = ~(_GEN_626 == _GEN_926) ? _GEN_1109 : grid_182; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1711 = ~(_GEN_626 == _GEN_926) ? _GEN_1110 : grid_183; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1712 = ~(_GEN_626 == _GEN_926) ? _GEN_1111 : grid_184; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1713 = ~(_GEN_626 == _GEN_926) ? _GEN_1112 : grid_185; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1714 = ~(_GEN_626 == _GEN_926) ? _GEN_1113 : grid_186; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1715 = ~(_GEN_626 == _GEN_926) ? _GEN_1114 : grid_187; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1716 = ~(_GEN_626 == _GEN_926) ? _GEN_1115 : grid_188; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1717 = ~(_GEN_626 == _GEN_926) ? _GEN_1116 : grid_189; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1718 = ~(_GEN_626 == _GEN_926) ? _GEN_1117 : grid_190; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1719 = ~(_GEN_626 == _GEN_926) ? _GEN_1118 : grid_191; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1720 = ~(_GEN_626 == _GEN_926) ? _GEN_1119 : grid_192; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1721 = ~(_GEN_626 == _GEN_926) ? _GEN_1120 : grid_193; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1722 = ~(_GEN_626 == _GEN_926) ? _GEN_1121 : grid_194; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1723 = ~(_GEN_626 == _GEN_926) ? _GEN_1122 : grid_195; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1724 = ~(_GEN_626 == _GEN_926) ? _GEN_1123 : grid_196; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1725 = ~(_GEN_626 == _GEN_926) ? _GEN_1124 : grid_197; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1726 = ~(_GEN_626 == _GEN_926) ? _GEN_1125 : grid_198; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1727 = ~(_GEN_626 == _GEN_926) ? _GEN_1126 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1728 = ~(_GEN_626 == _GEN_926) ? _GEN_1127 : grid_200; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1729 = ~(_GEN_626 == _GEN_926) ? _GEN_1128 : grid_201; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1730 = ~(_GEN_626 == _GEN_926) ? _GEN_1129 : grid_202; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1731 = ~(_GEN_626 == _GEN_926) ? _GEN_1130 : grid_203; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1732 = ~(_GEN_626 == _GEN_926) ? _GEN_1131 : grid_204; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1733 = ~(_GEN_626 == _GEN_926) ? _GEN_1132 : grid_205; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1734 = ~(_GEN_626 == _GEN_926) ? _GEN_1133 : grid_206; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1735 = ~(_GEN_626 == _GEN_926) ? _GEN_1134 : grid_207; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1736 = ~(_GEN_626 == _GEN_926) ? _GEN_1135 : grid_208; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1737 = ~(_GEN_626 == _GEN_926) ? _GEN_1136 : grid_209; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1738 = ~(_GEN_626 == _GEN_926) ? _GEN_1137 : grid_210; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1739 = ~(_GEN_626 == _GEN_926) ? _GEN_1138 : grid_211; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1740 = ~(_GEN_626 == _GEN_926) ? _GEN_1139 : grid_212; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1741 = ~(_GEN_626 == _GEN_926) ? _GEN_1140 : grid_213; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1742 = ~(_GEN_626 == _GEN_926) ? _GEN_1141 : grid_214; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1743 = ~(_GEN_626 == _GEN_926) ? _GEN_1142 : grid_215; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1744 = ~(_GEN_626 == _GEN_926) ? _GEN_1143 : grid_216; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1745 = ~(_GEN_626 == _GEN_926) ? _GEN_1144 : grid_217; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1746 = ~(_GEN_626 == _GEN_926) ? _GEN_1145 : grid_218; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1747 = ~(_GEN_626 == _GEN_926) ? _GEN_1146 : grid_219; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1748 = ~(_GEN_626 == _GEN_926) ? _GEN_1147 : grid_220; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1749 = ~(_GEN_626 == _GEN_926) ? _GEN_1148 : grid_221; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1750 = ~(_GEN_626 == _GEN_926) ? _GEN_1149 : grid_222; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1751 = ~(_GEN_626 == _GEN_926) ? _GEN_1150 : grid_223; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1752 = ~(_GEN_626 == _GEN_926) ? _GEN_1151 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1753 = ~(_GEN_626 == _GEN_926) ? _GEN_1152 : grid_225; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1754 = ~(_GEN_626 == _GEN_926) ? _GEN_1153 : grid_226; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1755 = ~(_GEN_626 == _GEN_926) ? _GEN_1154 : grid_227; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1756 = ~(_GEN_626 == _GEN_926) ? _GEN_1155 : grid_228; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1757 = ~(_GEN_626 == _GEN_926) ? _GEN_1156 : grid_229; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1758 = ~(_GEN_626 == _GEN_926) ? _GEN_1157 : grid_230; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1759 = ~(_GEN_626 == _GEN_926) ? _GEN_1158 : grid_231; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1760 = ~(_GEN_626 == _GEN_926) ? _GEN_1159 : grid_232; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1761 = ~(_GEN_626 == _GEN_926) ? _GEN_1160 : grid_233; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1762 = ~(_GEN_626 == _GEN_926) ? _GEN_1161 : grid_234; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1763 = ~(_GEN_626 == _GEN_926) ? _GEN_1162 : grid_235; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1764 = ~(_GEN_626 == _GEN_926) ? _GEN_1163 : grid_236; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1765 = ~(_GEN_626 == _GEN_926) ? _GEN_1164 : grid_237; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1766 = ~(_GEN_626 == _GEN_926) ? _GEN_1165 : grid_238; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1767 = ~(_GEN_626 == _GEN_926) ? _GEN_1166 : grid_239; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1768 = ~(_GEN_626 == _GEN_926) ? _GEN_1167 : grid_240; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1769 = ~(_GEN_626 == _GEN_926) ? _GEN_1168 : grid_241; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1770 = ~(_GEN_626 == _GEN_926) ? _GEN_1169 : grid_242; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1771 = ~(_GEN_626 == _GEN_926) ? _GEN_1170 : grid_243; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1772 = ~(_GEN_626 == _GEN_926) ? _GEN_1171 : grid_244; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1773 = ~(_GEN_626 == _GEN_926) ? _GEN_1172 : grid_245; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1774 = ~(_GEN_626 == _GEN_926) ? _GEN_1173 : grid_246; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1775 = ~(_GEN_626 == _GEN_926) ? _GEN_1174 : grid_247; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1776 = ~(_GEN_626 == _GEN_926) ? _GEN_1175 : grid_248; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1777 = ~(_GEN_626 == _GEN_926) ? _GEN_1176 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1778 = ~(_GEN_626 == _GEN_926) ? _GEN_1177 : grid_250; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1779 = ~(_GEN_626 == _GEN_926) ? _GEN_1178 : grid_251; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1780 = ~(_GEN_626 == _GEN_926) ? _GEN_1179 : grid_252; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1781 = ~(_GEN_626 == _GEN_926) ? _GEN_1180 : grid_253; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1782 = ~(_GEN_626 == _GEN_926) ? _GEN_1181 : grid_254; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1783 = ~(_GEN_626 == _GEN_926) ? _GEN_1182 : grid_255; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1784 = ~(_GEN_626 == _GEN_926) ? _GEN_1183 : grid_256; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1785 = ~(_GEN_626 == _GEN_926) ? _GEN_1184 : grid_257; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1786 = ~(_GEN_626 == _GEN_926) ? _GEN_1185 : grid_258; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1787 = ~(_GEN_626 == _GEN_926) ? _GEN_1186 : grid_259; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1788 = ~(_GEN_626 == _GEN_926) ? _GEN_1187 : grid_260; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1789 = ~(_GEN_626 == _GEN_926) ? _GEN_1188 : grid_261; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1790 = ~(_GEN_626 == _GEN_926) ? _GEN_1189 : grid_262; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1791 = ~(_GEN_626 == _GEN_926) ? _GEN_1190 : grid_263; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1792 = ~(_GEN_626 == _GEN_926) ? _GEN_1191 : grid_264; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1793 = ~(_GEN_626 == _GEN_926) ? _GEN_1192 : grid_265; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1794 = ~(_GEN_626 == _GEN_926) ? _GEN_1193 : grid_266; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1795 = ~(_GEN_626 == _GEN_926) ? _GEN_1194 : grid_267; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1796 = ~(_GEN_626 == _GEN_926) ? _GEN_1195 : grid_268; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1797 = ~(_GEN_626 == _GEN_926) ? _GEN_1196 : grid_269; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1798 = ~(_GEN_626 == _GEN_926) ? _GEN_1197 : grid_270; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1799 = ~(_GEN_626 == _GEN_926) ? _GEN_1198 : grid_271; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1800 = ~(_GEN_626 == _GEN_926) ? _GEN_1199 : grid_272; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1801 = ~(_GEN_626 == _GEN_926) ? _GEN_1200 : grid_273; // @[\\src\\main\\scala\\GameLogic.scala 230:53 88:21]
  wire [1:0] _GEN_1802 = ~(_GEN_626 == _GEN_926) ? _GEN_1201 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 91:23]
  wire [1:0] _GEN_1803 = ~(_GEN_626 == _GEN_926) ? _GEN_1202 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1804 = ~(_GEN_626 == _GEN_926) ? _GEN_1203 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1805 = ~(_GEN_626 == _GEN_926) ? _GEN_1204 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1806 = ~(_GEN_626 == _GEN_926) ? _GEN_1205 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1807 = ~(_GEN_626 == _GEN_926) ? _GEN_1206 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1808 = ~(_GEN_626 == _GEN_926) ? _GEN_1207 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1809 = ~(_GEN_626 == _GEN_926) ? _GEN_1208 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1810 = ~(_GEN_626 == _GEN_926) ? _GEN_1209 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1811 = ~(_GEN_626 == _GEN_926) ? _GEN_1210 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1812 = ~(_GEN_626 == _GEN_926) ? _GEN_1211 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1813 = ~(_GEN_626 == _GEN_926) ? _GEN_1212 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1814 = ~(_GEN_626 == _GEN_926) ? _GEN_1213 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1815 = ~(_GEN_626 == _GEN_926) ? _GEN_1214 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1816 = ~(_GEN_626 == _GEN_926) ? _GEN_1215 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1817 = ~(_GEN_626 == _GEN_926) ? _GEN_1216 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1818 = ~(_GEN_626 == _GEN_926) ? _GEN_1217 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1819 = ~(_GEN_626 == _GEN_926) ? _GEN_1218 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1820 = ~(_GEN_626 == _GEN_926) ? _GEN_1219 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1821 = ~(_GEN_626 == _GEN_926) ? _GEN_1220 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1822 = ~(_GEN_626 == _GEN_926) ? _GEN_1221 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1823 = ~(_GEN_626 == _GEN_926) ? _GEN_1222 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1824 = ~(_GEN_626 == _GEN_926) ? _GEN_1223 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1825 = ~(_GEN_626 == _GEN_926) ? _GEN_1224 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1826 = ~(_GEN_626 == _GEN_926) ? _GEN_1225 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [1:0] _GEN_1827 = ~(_GEN_626 == _GEN_926) ? _GEN_1226 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 230:53 96:21]
  wire [3:0] _currentBlock_T_1 = currentBlock + 4'h1; // @[\\src\\main\\scala\\GameLogic.scala 234:42]
  wire [1:0] _GEN_1828 = currentBlock == 4'h9 ? 2'h3 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 220:41 221:22 137:25]
  wire [3:0] _GEN_1829 = currentBlock == 4'h9 ? 4'h0 : _currentBlock_T_1; // @[\\src\\main\\scala\\GameLogic.scala 220:41 222:26 234:26]
  wire [8:0] _GEN_1830 = currentBlock == 4'h9 ? 9'h0 : index; // @[\\src\\main\\scala\\GameLogic.scala 129:29 220:41 228:39]
  wire [4:0] _GEN_1831 = currentBlock == 4'h9 ? 5'h0 : _GEN_1527; // @[\\src\\main\\scala\\GameLogic.scala 128:26 220:41]
  wire [1:0] _GEN_1832 = currentBlock == 4'h9 ? 2'h1 : _GEN_1528; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1833 = currentBlock == 4'h9 ? 2'h1 : _GEN_1529; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1834 = currentBlock == 4'h9 ? 2'h1 : _GEN_1530; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1835 = currentBlock == 4'h9 ? 2'h1 : _GEN_1531; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1836 = currentBlock == 4'h9 ? 2'h1 : _GEN_1532; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1837 = currentBlock == 4'h9 ? 2'h1 : _GEN_1533; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1838 = currentBlock == 4'h9 ? 2'h1 : _GEN_1534; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1839 = currentBlock == 4'h9 ? 2'h1 : _GEN_1535; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1840 = currentBlock == 4'h9 ? 2'h1 : _GEN_1536; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1841 = currentBlock == 4'h9 ? 2'h1 : _GEN_1537; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1842 = currentBlock == 4'h9 ? 2'h1 : _GEN_1538; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1843 = currentBlock == 4'h9 ? 2'h1 : _GEN_1539; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1844 = currentBlock == 4'h9 ? 2'h1 : _GEN_1540; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1845 = currentBlock == 4'h9 ? 2'h1 : _GEN_1541; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1846 = currentBlock == 4'h9 ? 2'h1 : _GEN_1542; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1847 = currentBlock == 4'h9 ? 2'h1 : _GEN_1543; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1848 = currentBlock == 4'h9 ? 2'h1 : _GEN_1544; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1849 = currentBlock == 4'h9 ? 2'h1 : _GEN_1545; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1850 = currentBlock == 4'h9 ? 2'h1 : _GEN_1546; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1851 = currentBlock == 4'h9 ? 2'h1 : _GEN_1547; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1852 = currentBlock == 4'h9 ? 2'h1 : _GEN_1548; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1853 = currentBlock == 4'h9 ? 2'h1 : _GEN_1549; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1854 = currentBlock == 4'h9 ? 2'h1 : _GEN_1550; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1855 = currentBlock == 4'h9 ? 2'h1 : _GEN_1551; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1856 = currentBlock == 4'h9 ? 2'h1 : _GEN_1552; // @[\\src\\main\\scala\\GameLogic.scala 220:41 95:13]
  wire [1:0] _GEN_1857 = currentBlock == 4'h9 ? grid_25 : _GEN_1553; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1858 = currentBlock == 4'h9 ? grid_26 : _GEN_1554; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1859 = currentBlock == 4'h9 ? grid_27 : _GEN_1555; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1860 = currentBlock == 4'h9 ? grid_28 : _GEN_1556; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1861 = currentBlock == 4'h9 ? grid_29 : _GEN_1557; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1862 = currentBlock == 4'h9 ? grid_30 : _GEN_1558; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1863 = currentBlock == 4'h9 ? grid_31 : _GEN_1559; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1864 = currentBlock == 4'h9 ? grid_32 : _GEN_1560; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1865 = currentBlock == 4'h9 ? grid_33 : _GEN_1561; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1866 = currentBlock == 4'h9 ? grid_34 : _GEN_1562; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1867 = currentBlock == 4'h9 ? grid_35 : _GEN_1563; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1868 = currentBlock == 4'h9 ? grid_36 : _GEN_1564; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1869 = currentBlock == 4'h9 ? grid_37 : _GEN_1565; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1870 = currentBlock == 4'h9 ? grid_38 : _GEN_1566; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1871 = currentBlock == 4'h9 ? grid_39 : _GEN_1567; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1872 = currentBlock == 4'h9 ? grid_40 : _GEN_1568; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1873 = currentBlock == 4'h9 ? grid_41 : _GEN_1569; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1874 = currentBlock == 4'h9 ? grid_42 : _GEN_1570; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1875 = currentBlock == 4'h9 ? grid_43 : _GEN_1571; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1876 = currentBlock == 4'h9 ? grid_44 : _GEN_1572; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1877 = currentBlock == 4'h9 ? grid_45 : _GEN_1573; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1878 = currentBlock == 4'h9 ? grid_46 : _GEN_1574; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1879 = currentBlock == 4'h9 ? grid_47 : _GEN_1575; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1880 = currentBlock == 4'h9 ? grid_48 : _GEN_1576; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1881 = currentBlock == 4'h9 ? 2'h1 : _GEN_1577; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_1882 = currentBlock == 4'h9 ? grid_50 : _GEN_1578; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1883 = currentBlock == 4'h9 ? grid_51 : _GEN_1579; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1884 = currentBlock == 4'h9 ? grid_52 : _GEN_1580; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1885 = currentBlock == 4'h9 ? grid_53 : _GEN_1581; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1886 = currentBlock == 4'h9 ? grid_54 : _GEN_1582; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1887 = currentBlock == 4'h9 ? grid_55 : _GEN_1583; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1888 = currentBlock == 4'h9 ? grid_56 : _GEN_1584; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1889 = currentBlock == 4'h9 ? grid_57 : _GEN_1585; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1890 = currentBlock == 4'h9 ? grid_58 : _GEN_1586; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1891 = currentBlock == 4'h9 ? grid_59 : _GEN_1587; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1892 = currentBlock == 4'h9 ? grid_60 : _GEN_1588; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1893 = currentBlock == 4'h9 ? grid_61 : _GEN_1589; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1894 = currentBlock == 4'h9 ? grid_62 : _GEN_1590; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1895 = currentBlock == 4'h9 ? grid_63 : _GEN_1591; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1896 = currentBlock == 4'h9 ? grid_64 : _GEN_1592; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1897 = currentBlock == 4'h9 ? grid_65 : _GEN_1593; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1898 = currentBlock == 4'h9 ? grid_66 : _GEN_1594; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1899 = currentBlock == 4'h9 ? grid_67 : _GEN_1595; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1900 = currentBlock == 4'h9 ? grid_68 : _GEN_1596; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1901 = currentBlock == 4'h9 ? grid_69 : _GEN_1597; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1902 = currentBlock == 4'h9 ? grid_70 : _GEN_1598; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1903 = currentBlock == 4'h9 ? grid_71 : _GEN_1599; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1904 = currentBlock == 4'h9 ? grid_72 : _GEN_1600; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1905 = currentBlock == 4'h9 ? grid_73 : _GEN_1601; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1906 = currentBlock == 4'h9 ? 2'h1 : _GEN_1602; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_1907 = currentBlock == 4'h9 ? grid_75 : _GEN_1603; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1908 = currentBlock == 4'h9 ? grid_76 : _GEN_1604; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1909 = currentBlock == 4'h9 ? grid_77 : _GEN_1605; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1910 = currentBlock == 4'h9 ? grid_78 : _GEN_1606; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1911 = currentBlock == 4'h9 ? grid_79 : _GEN_1607; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1912 = currentBlock == 4'h9 ? grid_80 : _GEN_1608; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1913 = currentBlock == 4'h9 ? grid_81 : _GEN_1609; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1914 = currentBlock == 4'h9 ? grid_82 : _GEN_1610; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1915 = currentBlock == 4'h9 ? grid_83 : _GEN_1611; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1916 = currentBlock == 4'h9 ? grid_84 : _GEN_1612; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1917 = currentBlock == 4'h9 ? grid_85 : _GEN_1613; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1918 = currentBlock == 4'h9 ? grid_86 : _GEN_1614; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1919 = currentBlock == 4'h9 ? grid_87 : _GEN_1615; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1920 = currentBlock == 4'h9 ? grid_88 : _GEN_1616; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1921 = currentBlock == 4'h9 ? grid_89 : _GEN_1617; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1922 = currentBlock == 4'h9 ? grid_90 : _GEN_1618; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1923 = currentBlock == 4'h9 ? grid_91 : _GEN_1619; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1924 = currentBlock == 4'h9 ? grid_92 : _GEN_1620; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1925 = currentBlock == 4'h9 ? grid_93 : _GEN_1621; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1926 = currentBlock == 4'h9 ? grid_94 : _GEN_1622; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1927 = currentBlock == 4'h9 ? grid_95 : _GEN_1623; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1928 = currentBlock == 4'h9 ? grid_96 : _GEN_1624; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1929 = currentBlock == 4'h9 ? grid_97 : _GEN_1625; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1930 = currentBlock == 4'h9 ? grid_98 : _GEN_1626; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1931 = currentBlock == 4'h9 ? 2'h1 : _GEN_1627; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_1932 = currentBlock == 4'h9 ? grid_100 : _GEN_1628; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1933 = currentBlock == 4'h9 ? grid_101 : _GEN_1629; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1934 = currentBlock == 4'h9 ? grid_102 : _GEN_1630; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1935 = currentBlock == 4'h9 ? grid_103 : _GEN_1631; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1936 = currentBlock == 4'h9 ? grid_104 : _GEN_1632; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1937 = currentBlock == 4'h9 ? grid_105 : _GEN_1633; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1938 = currentBlock == 4'h9 ? grid_106 : _GEN_1634; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1939 = currentBlock == 4'h9 ? grid_107 : _GEN_1635; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1940 = currentBlock == 4'h9 ? grid_108 : _GEN_1636; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1941 = currentBlock == 4'h9 ? grid_109 : _GEN_1637; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1942 = currentBlock == 4'h9 ? grid_110 : _GEN_1638; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1943 = currentBlock == 4'h9 ? grid_111 : _GEN_1639; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1944 = currentBlock == 4'h9 ? grid_112 : _GEN_1640; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1945 = currentBlock == 4'h9 ? grid_113 : _GEN_1641; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1946 = currentBlock == 4'h9 ? grid_114 : _GEN_1642; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1947 = currentBlock == 4'h9 ? grid_115 : _GEN_1643; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1948 = currentBlock == 4'h9 ? grid_116 : _GEN_1644; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1949 = currentBlock == 4'h9 ? grid_117 : _GEN_1645; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1950 = currentBlock == 4'h9 ? grid_118 : _GEN_1646; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1951 = currentBlock == 4'h9 ? grid_119 : _GEN_1647; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1952 = currentBlock == 4'h9 ? grid_120 : _GEN_1648; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1953 = currentBlock == 4'h9 ? grid_121 : _GEN_1649; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1954 = currentBlock == 4'h9 ? grid_122 : _GEN_1650; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1955 = currentBlock == 4'h9 ? grid_123 : _GEN_1651; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1956 = currentBlock == 4'h9 ? 2'h1 : _GEN_1652; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_1957 = currentBlock == 4'h9 ? grid_125 : _GEN_1653; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1958 = currentBlock == 4'h9 ? grid_126 : _GEN_1654; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1959 = currentBlock == 4'h9 ? grid_127 : _GEN_1655; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1960 = currentBlock == 4'h9 ? grid_128 : _GEN_1656; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1961 = currentBlock == 4'h9 ? grid_129 : _GEN_1657; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1962 = currentBlock == 4'h9 ? grid_130 : _GEN_1658; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1963 = currentBlock == 4'h9 ? grid_131 : _GEN_1659; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1964 = currentBlock == 4'h9 ? grid_132 : _GEN_1660; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1965 = currentBlock == 4'h9 ? grid_133 : _GEN_1661; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1966 = currentBlock == 4'h9 ? grid_134 : _GEN_1662; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1967 = currentBlock == 4'h9 ? grid_135 : _GEN_1663; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1968 = currentBlock == 4'h9 ? grid_136 : _GEN_1664; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1969 = currentBlock == 4'h9 ? grid_137 : _GEN_1665; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1970 = currentBlock == 4'h9 ? grid_138 : _GEN_1666; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1971 = currentBlock == 4'h9 ? grid_139 : _GEN_1667; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1972 = currentBlock == 4'h9 ? grid_140 : _GEN_1668; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1973 = currentBlock == 4'h9 ? grid_141 : _GEN_1669; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1974 = currentBlock == 4'h9 ? grid_142 : _GEN_1670; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1975 = currentBlock == 4'h9 ? grid_143 : _GEN_1671; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1976 = currentBlock == 4'h9 ? grid_144 : _GEN_1672; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1977 = currentBlock == 4'h9 ? grid_145 : _GEN_1673; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1978 = currentBlock == 4'h9 ? grid_146 : _GEN_1674; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1979 = currentBlock == 4'h9 ? grid_147 : _GEN_1675; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1980 = currentBlock == 4'h9 ? grid_148 : _GEN_1676; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1981 = currentBlock == 4'h9 ? 2'h1 : _GEN_1677; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_1982 = currentBlock == 4'h9 ? grid_150 : _GEN_1678; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1983 = currentBlock == 4'h9 ? grid_151 : _GEN_1679; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1984 = currentBlock == 4'h9 ? grid_152 : _GEN_1680; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1985 = currentBlock == 4'h9 ? grid_153 : _GEN_1681; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1986 = currentBlock == 4'h9 ? grid_154 : _GEN_1682; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1987 = currentBlock == 4'h9 ? grid_155 : _GEN_1683; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1988 = currentBlock == 4'h9 ? grid_156 : _GEN_1684; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1989 = currentBlock == 4'h9 ? grid_157 : _GEN_1685; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1990 = currentBlock == 4'h9 ? grid_158 : _GEN_1686; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1991 = currentBlock == 4'h9 ? grid_159 : _GEN_1687; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1992 = currentBlock == 4'h9 ? grid_160 : _GEN_1688; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1993 = currentBlock == 4'h9 ? grid_161 : _GEN_1689; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1994 = currentBlock == 4'h9 ? grid_162 : _GEN_1690; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1995 = currentBlock == 4'h9 ? grid_163 : _GEN_1691; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1996 = currentBlock == 4'h9 ? grid_164 : _GEN_1692; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1997 = currentBlock == 4'h9 ? grid_165 : _GEN_1693; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1998 = currentBlock == 4'h9 ? grid_166 : _GEN_1694; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_1999 = currentBlock == 4'h9 ? grid_167 : _GEN_1695; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2000 = currentBlock == 4'h9 ? grid_168 : _GEN_1696; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2001 = currentBlock == 4'h9 ? grid_169 : _GEN_1697; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2002 = currentBlock == 4'h9 ? grid_170 : _GEN_1698; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2003 = currentBlock == 4'h9 ? grid_171 : _GEN_1699; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2004 = currentBlock == 4'h9 ? grid_172 : _GEN_1700; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2005 = currentBlock == 4'h9 ? grid_173 : _GEN_1701; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2006 = currentBlock == 4'h9 ? 2'h1 : _GEN_1702; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_2007 = currentBlock == 4'h9 ? grid_175 : _GEN_1703; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2008 = currentBlock == 4'h9 ? grid_176 : _GEN_1704; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2009 = currentBlock == 4'h9 ? grid_177 : _GEN_1705; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2010 = currentBlock == 4'h9 ? grid_178 : _GEN_1706; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2011 = currentBlock == 4'h9 ? grid_179 : _GEN_1707; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2012 = currentBlock == 4'h9 ? grid_180 : _GEN_1708; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2013 = currentBlock == 4'h9 ? grid_181 : _GEN_1709; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2014 = currentBlock == 4'h9 ? grid_182 : _GEN_1710; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2015 = currentBlock == 4'h9 ? grid_183 : _GEN_1711; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2016 = currentBlock == 4'h9 ? grid_184 : _GEN_1712; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2017 = currentBlock == 4'h9 ? grid_185 : _GEN_1713; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2018 = currentBlock == 4'h9 ? grid_186 : _GEN_1714; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2019 = currentBlock == 4'h9 ? grid_187 : _GEN_1715; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2020 = currentBlock == 4'h9 ? grid_188 : _GEN_1716; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2021 = currentBlock == 4'h9 ? grid_189 : _GEN_1717; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2022 = currentBlock == 4'h9 ? grid_190 : _GEN_1718; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2023 = currentBlock == 4'h9 ? grid_191 : _GEN_1719; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2024 = currentBlock == 4'h9 ? grid_192 : _GEN_1720; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2025 = currentBlock == 4'h9 ? grid_193 : _GEN_1721; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2026 = currentBlock == 4'h9 ? grid_194 : _GEN_1722; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2027 = currentBlock == 4'h9 ? grid_195 : _GEN_1723; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2028 = currentBlock == 4'h9 ? grid_196 : _GEN_1724; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2029 = currentBlock == 4'h9 ? grid_197 : _GEN_1725; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2030 = currentBlock == 4'h9 ? grid_198 : _GEN_1726; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2031 = currentBlock == 4'h9 ? 2'h1 : _GEN_1727; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_2032 = currentBlock == 4'h9 ? grid_200 : _GEN_1728; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2033 = currentBlock == 4'h9 ? grid_201 : _GEN_1729; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2034 = currentBlock == 4'h9 ? grid_202 : _GEN_1730; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2035 = currentBlock == 4'h9 ? grid_203 : _GEN_1731; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2036 = currentBlock == 4'h9 ? grid_204 : _GEN_1732; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2037 = currentBlock == 4'h9 ? grid_205 : _GEN_1733; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2038 = currentBlock == 4'h9 ? grid_206 : _GEN_1734; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2039 = currentBlock == 4'h9 ? grid_207 : _GEN_1735; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2040 = currentBlock == 4'h9 ? grid_208 : _GEN_1736; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2041 = currentBlock == 4'h9 ? grid_209 : _GEN_1737; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2042 = currentBlock == 4'h9 ? grid_210 : _GEN_1738; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2043 = currentBlock == 4'h9 ? grid_211 : _GEN_1739; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2044 = currentBlock == 4'h9 ? grid_212 : _GEN_1740; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2045 = currentBlock == 4'h9 ? grid_213 : _GEN_1741; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2046 = currentBlock == 4'h9 ? grid_214 : _GEN_1742; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2047 = currentBlock == 4'h9 ? grid_215 : _GEN_1743; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2048 = currentBlock == 4'h9 ? grid_216 : _GEN_1744; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2049 = currentBlock == 4'h9 ? grid_217 : _GEN_1745; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2050 = currentBlock == 4'h9 ? grid_218 : _GEN_1746; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2051 = currentBlock == 4'h9 ? grid_219 : _GEN_1747; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2052 = currentBlock == 4'h9 ? grid_220 : _GEN_1748; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2053 = currentBlock == 4'h9 ? grid_221 : _GEN_1749; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2054 = currentBlock == 4'h9 ? grid_222 : _GEN_1750; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2055 = currentBlock == 4'h9 ? grid_223 : _GEN_1751; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2056 = currentBlock == 4'h9 ? 2'h1 : _GEN_1752; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_2057 = currentBlock == 4'h9 ? grid_225 : _GEN_1753; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2058 = currentBlock == 4'h9 ? grid_226 : _GEN_1754; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2059 = currentBlock == 4'h9 ? grid_227 : _GEN_1755; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2060 = currentBlock == 4'h9 ? grid_228 : _GEN_1756; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2061 = currentBlock == 4'h9 ? grid_229 : _GEN_1757; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2062 = currentBlock == 4'h9 ? grid_230 : _GEN_1758; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2063 = currentBlock == 4'h9 ? grid_231 : _GEN_1759; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2064 = currentBlock == 4'h9 ? grid_232 : _GEN_1760; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2065 = currentBlock == 4'h9 ? grid_233 : _GEN_1761; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2066 = currentBlock == 4'h9 ? grid_234 : _GEN_1762; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2067 = currentBlock == 4'h9 ? grid_235 : _GEN_1763; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2068 = currentBlock == 4'h9 ? grid_236 : _GEN_1764; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2069 = currentBlock == 4'h9 ? grid_237 : _GEN_1765; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2070 = currentBlock == 4'h9 ? grid_238 : _GEN_1766; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2071 = currentBlock == 4'h9 ? grid_239 : _GEN_1767; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2072 = currentBlock == 4'h9 ? grid_240 : _GEN_1768; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2073 = currentBlock == 4'h9 ? grid_241 : _GEN_1769; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2074 = currentBlock == 4'h9 ? grid_242 : _GEN_1770; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2075 = currentBlock == 4'h9 ? grid_243 : _GEN_1771; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2076 = currentBlock == 4'h9 ? grid_244 : _GEN_1772; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2077 = currentBlock == 4'h9 ? grid_245 : _GEN_1773; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2078 = currentBlock == 4'h9 ? grid_246 : _GEN_1774; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2079 = currentBlock == 4'h9 ? grid_247 : _GEN_1775; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2080 = currentBlock == 4'h9 ? grid_248 : _GEN_1776; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2081 = currentBlock == 4'h9 ? 2'h1 : _GEN_1777; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_2082 = currentBlock == 4'h9 ? grid_250 : _GEN_1778; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2083 = currentBlock == 4'h9 ? grid_251 : _GEN_1779; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2084 = currentBlock == 4'h9 ? grid_252 : _GEN_1780; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2085 = currentBlock == 4'h9 ? grid_253 : _GEN_1781; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2086 = currentBlock == 4'h9 ? grid_254 : _GEN_1782; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2087 = currentBlock == 4'h9 ? grid_255 : _GEN_1783; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2088 = currentBlock == 4'h9 ? grid_256 : _GEN_1784; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2089 = currentBlock == 4'h9 ? grid_257 : _GEN_1785; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2090 = currentBlock == 4'h9 ? grid_258 : _GEN_1786; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2091 = currentBlock == 4'h9 ? grid_259 : _GEN_1787; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2092 = currentBlock == 4'h9 ? grid_260 : _GEN_1788; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2093 = currentBlock == 4'h9 ? grid_261 : _GEN_1789; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2094 = currentBlock == 4'h9 ? grid_262 : _GEN_1790; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2095 = currentBlock == 4'h9 ? grid_263 : _GEN_1791; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2096 = currentBlock == 4'h9 ? grid_264 : _GEN_1792; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2097 = currentBlock == 4'h9 ? grid_265 : _GEN_1793; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2098 = currentBlock == 4'h9 ? grid_266 : _GEN_1794; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2099 = currentBlock == 4'h9 ? grid_267 : _GEN_1795; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2100 = currentBlock == 4'h9 ? grid_268 : _GEN_1796; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2101 = currentBlock == 4'h9 ? grid_269 : _GEN_1797; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2102 = currentBlock == 4'h9 ? grid_270 : _GEN_1798; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2103 = currentBlock == 4'h9 ? grid_271 : _GEN_1799; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2104 = currentBlock == 4'h9 ? grid_272 : _GEN_1800; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2105 = currentBlock == 4'h9 ? grid_273 : _GEN_1801; // @[\\src\\main\\scala\\GameLogic.scala 220:41 88:21]
  wire [1:0] _GEN_2106 = currentBlock == 4'h9 ? 2'h1 : _GEN_1802; // @[\\src\\main\\scala\\GameLogic.scala 220:41 91:23]
  wire [1:0] _GEN_2107 = currentBlock == 4'h9 ? 2'h1 : _GEN_1803; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2108 = currentBlock == 4'h9 ? 2'h1 : _GEN_1804; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2109 = currentBlock == 4'h9 ? 2'h1 : _GEN_1805; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2110 = currentBlock == 4'h9 ? 2'h1 : _GEN_1806; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2111 = currentBlock == 4'h9 ? 2'h1 : _GEN_1807; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2112 = currentBlock == 4'h9 ? 2'h1 : _GEN_1808; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2113 = currentBlock == 4'h9 ? 2'h1 : _GEN_1809; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2114 = currentBlock == 4'h9 ? 2'h1 : _GEN_1810; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2115 = currentBlock == 4'h9 ? 2'h1 : _GEN_1811; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2116 = currentBlock == 4'h9 ? 2'h1 : _GEN_1812; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2117 = currentBlock == 4'h9 ? 2'h1 : _GEN_1813; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2118 = currentBlock == 4'h9 ? 2'h1 : _GEN_1814; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2119 = currentBlock == 4'h9 ? 2'h1 : _GEN_1815; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2120 = currentBlock == 4'h9 ? 2'h1 : _GEN_1816; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2121 = currentBlock == 4'h9 ? 2'h1 : _GEN_1817; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2122 = currentBlock == 4'h9 ? 2'h1 : _GEN_1818; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2123 = currentBlock == 4'h9 ? 2'h1 : _GEN_1819; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2124 = currentBlock == 4'h9 ? 2'h1 : _GEN_1820; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2125 = currentBlock == 4'h9 ? 2'h1 : _GEN_1821; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2126 = currentBlock == 4'h9 ? 2'h1 : _GEN_1822; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2127 = currentBlock == 4'h9 ? 2'h1 : _GEN_1823; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2128 = currentBlock == 4'h9 ? 2'h1 : _GEN_1824; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2129 = currentBlock == 4'h9 ? 2'h1 : _GEN_1825; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2130 = currentBlock == 4'h9 ? 2'h1 : _GEN_1826; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2131 = currentBlock == 4'h9 ? 2'h1 : _GEN_1827; // @[\\src\\main\\scala\\GameLogic.scala 220:41 96:21]
  wire [1:0] _GEN_2132 = 2'h2 == currentTask ? _GEN_1828 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 137:25 196:27]
  wire [3:0] _GEN_2133 = 2'h2 == currentTask ? _GEN_1829 : currentBlock; // @[\\src\\main\\scala\\GameLogic.scala 196:27 84:29]
  wire [8:0] _GEN_2134 = 2'h2 == currentTask ? _GEN_1830 : 9'h0; // @[\\src\\main\\scala\\GameLogic.scala 196:27 129:29]
  wire [4:0] _GEN_2135 = 2'h2 == currentTask ? _GEN_1831 : 5'h0; // @[\\src\\main\\scala\\GameLogic.scala 128:26 196:27]
  wire [1:0] _GEN_2136 = 2'h2 == currentTask ? _GEN_1832 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2137 = 2'h2 == currentTask ? _GEN_1833 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2138 = 2'h2 == currentTask ? _GEN_1834 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2139 = 2'h2 == currentTask ? _GEN_1835 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2140 = 2'h2 == currentTask ? _GEN_1836 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2141 = 2'h2 == currentTask ? _GEN_1837 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2142 = 2'h2 == currentTask ? _GEN_1838 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2143 = 2'h2 == currentTask ? _GEN_1839 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2144 = 2'h2 == currentTask ? _GEN_1840 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2145 = 2'h2 == currentTask ? _GEN_1841 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2146 = 2'h2 == currentTask ? _GEN_1842 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2147 = 2'h2 == currentTask ? _GEN_1843 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2148 = 2'h2 == currentTask ? _GEN_1844 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2149 = 2'h2 == currentTask ? _GEN_1845 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2150 = 2'h2 == currentTask ? _GEN_1846 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2151 = 2'h2 == currentTask ? _GEN_1847 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2152 = 2'h2 == currentTask ? _GEN_1848 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2153 = 2'h2 == currentTask ? _GEN_1849 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2154 = 2'h2 == currentTask ? _GEN_1850 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2155 = 2'h2 == currentTask ? _GEN_1851 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2156 = 2'h2 == currentTask ? _GEN_1852 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2157 = 2'h2 == currentTask ? _GEN_1853 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2158 = 2'h2 == currentTask ? _GEN_1854 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2159 = 2'h2 == currentTask ? _GEN_1855 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2160 = 2'h2 == currentTask ? _GEN_1856 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 95:13]
  wire [1:0] _GEN_2161 = 2'h2 == currentTask ? _GEN_1857 : grid_25; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2162 = 2'h2 == currentTask ? _GEN_1858 : grid_26; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2163 = 2'h2 == currentTask ? _GEN_1859 : grid_27; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2164 = 2'h2 == currentTask ? _GEN_1860 : grid_28; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2165 = 2'h2 == currentTask ? _GEN_1861 : grid_29; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2166 = 2'h2 == currentTask ? _GEN_1862 : grid_30; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2167 = 2'h2 == currentTask ? _GEN_1863 : grid_31; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2168 = 2'h2 == currentTask ? _GEN_1864 : grid_32; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2169 = 2'h2 == currentTask ? _GEN_1865 : grid_33; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2170 = 2'h2 == currentTask ? _GEN_1866 : grid_34; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2171 = 2'h2 == currentTask ? _GEN_1867 : grid_35; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2172 = 2'h2 == currentTask ? _GEN_1868 : grid_36; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2173 = 2'h2 == currentTask ? _GEN_1869 : grid_37; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2174 = 2'h2 == currentTask ? _GEN_1870 : grid_38; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2175 = 2'h2 == currentTask ? _GEN_1871 : grid_39; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2176 = 2'h2 == currentTask ? _GEN_1872 : grid_40; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2177 = 2'h2 == currentTask ? _GEN_1873 : grid_41; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2178 = 2'h2 == currentTask ? _GEN_1874 : grid_42; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2179 = 2'h2 == currentTask ? _GEN_1875 : grid_43; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2180 = 2'h2 == currentTask ? _GEN_1876 : grid_44; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2181 = 2'h2 == currentTask ? _GEN_1877 : grid_45; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2182 = 2'h2 == currentTask ? _GEN_1878 : grid_46; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2183 = 2'h2 == currentTask ? _GEN_1879 : grid_47; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2184 = 2'h2 == currentTask ? _GEN_1880 : grid_48; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2185 = 2'h2 == currentTask ? _GEN_1881 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2186 = 2'h2 == currentTask ? _GEN_1882 : grid_50; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2187 = 2'h2 == currentTask ? _GEN_1883 : grid_51; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2188 = 2'h2 == currentTask ? _GEN_1884 : grid_52; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2189 = 2'h2 == currentTask ? _GEN_1885 : grid_53; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2190 = 2'h2 == currentTask ? _GEN_1886 : grid_54; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2191 = 2'h2 == currentTask ? _GEN_1887 : grid_55; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2192 = 2'h2 == currentTask ? _GEN_1888 : grid_56; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2193 = 2'h2 == currentTask ? _GEN_1889 : grid_57; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2194 = 2'h2 == currentTask ? _GEN_1890 : grid_58; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2195 = 2'h2 == currentTask ? _GEN_1891 : grid_59; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2196 = 2'h2 == currentTask ? _GEN_1892 : grid_60; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2197 = 2'h2 == currentTask ? _GEN_1893 : grid_61; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2198 = 2'h2 == currentTask ? _GEN_1894 : grid_62; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2199 = 2'h2 == currentTask ? _GEN_1895 : grid_63; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2200 = 2'h2 == currentTask ? _GEN_1896 : grid_64; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2201 = 2'h2 == currentTask ? _GEN_1897 : grid_65; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2202 = 2'h2 == currentTask ? _GEN_1898 : grid_66; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2203 = 2'h2 == currentTask ? _GEN_1899 : grid_67; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2204 = 2'h2 == currentTask ? _GEN_1900 : grid_68; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2205 = 2'h2 == currentTask ? _GEN_1901 : grid_69; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2206 = 2'h2 == currentTask ? _GEN_1902 : grid_70; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2207 = 2'h2 == currentTask ? _GEN_1903 : grid_71; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2208 = 2'h2 == currentTask ? _GEN_1904 : grid_72; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2209 = 2'h2 == currentTask ? _GEN_1905 : grid_73; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2210 = 2'h2 == currentTask ? _GEN_1906 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2211 = 2'h2 == currentTask ? _GEN_1907 : grid_75; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2212 = 2'h2 == currentTask ? _GEN_1908 : grid_76; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2213 = 2'h2 == currentTask ? _GEN_1909 : grid_77; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2214 = 2'h2 == currentTask ? _GEN_1910 : grid_78; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2215 = 2'h2 == currentTask ? _GEN_1911 : grid_79; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2216 = 2'h2 == currentTask ? _GEN_1912 : grid_80; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2217 = 2'h2 == currentTask ? _GEN_1913 : grid_81; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2218 = 2'h2 == currentTask ? _GEN_1914 : grid_82; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2219 = 2'h2 == currentTask ? _GEN_1915 : grid_83; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2220 = 2'h2 == currentTask ? _GEN_1916 : grid_84; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2221 = 2'h2 == currentTask ? _GEN_1917 : grid_85; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2222 = 2'h2 == currentTask ? _GEN_1918 : grid_86; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2223 = 2'h2 == currentTask ? _GEN_1919 : grid_87; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2224 = 2'h2 == currentTask ? _GEN_1920 : grid_88; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2225 = 2'h2 == currentTask ? _GEN_1921 : grid_89; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2226 = 2'h2 == currentTask ? _GEN_1922 : grid_90; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2227 = 2'h2 == currentTask ? _GEN_1923 : grid_91; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2228 = 2'h2 == currentTask ? _GEN_1924 : grid_92; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2229 = 2'h2 == currentTask ? _GEN_1925 : grid_93; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2230 = 2'h2 == currentTask ? _GEN_1926 : grid_94; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2231 = 2'h2 == currentTask ? _GEN_1927 : grid_95; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2232 = 2'h2 == currentTask ? _GEN_1928 : grid_96; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2233 = 2'h2 == currentTask ? _GEN_1929 : grid_97; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2234 = 2'h2 == currentTask ? _GEN_1930 : grid_98; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2235 = 2'h2 == currentTask ? _GEN_1931 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2236 = 2'h2 == currentTask ? _GEN_1932 : grid_100; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2237 = 2'h2 == currentTask ? _GEN_1933 : grid_101; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2238 = 2'h2 == currentTask ? _GEN_1934 : grid_102; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2239 = 2'h2 == currentTask ? _GEN_1935 : grid_103; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2240 = 2'h2 == currentTask ? _GEN_1936 : grid_104; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2241 = 2'h2 == currentTask ? _GEN_1937 : grid_105; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2242 = 2'h2 == currentTask ? _GEN_1938 : grid_106; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2243 = 2'h2 == currentTask ? _GEN_1939 : grid_107; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2244 = 2'h2 == currentTask ? _GEN_1940 : grid_108; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2245 = 2'h2 == currentTask ? _GEN_1941 : grid_109; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2246 = 2'h2 == currentTask ? _GEN_1942 : grid_110; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2247 = 2'h2 == currentTask ? _GEN_1943 : grid_111; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2248 = 2'h2 == currentTask ? _GEN_1944 : grid_112; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2249 = 2'h2 == currentTask ? _GEN_1945 : grid_113; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2250 = 2'h2 == currentTask ? _GEN_1946 : grid_114; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2251 = 2'h2 == currentTask ? _GEN_1947 : grid_115; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2252 = 2'h2 == currentTask ? _GEN_1948 : grid_116; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2253 = 2'h2 == currentTask ? _GEN_1949 : grid_117; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2254 = 2'h2 == currentTask ? _GEN_1950 : grid_118; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2255 = 2'h2 == currentTask ? _GEN_1951 : grid_119; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2256 = 2'h2 == currentTask ? _GEN_1952 : grid_120; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2257 = 2'h2 == currentTask ? _GEN_1953 : grid_121; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2258 = 2'h2 == currentTask ? _GEN_1954 : grid_122; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2259 = 2'h2 == currentTask ? _GEN_1955 : grid_123; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2260 = 2'h2 == currentTask ? _GEN_1956 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2261 = 2'h2 == currentTask ? _GEN_1957 : grid_125; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2262 = 2'h2 == currentTask ? _GEN_1958 : grid_126; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2263 = 2'h2 == currentTask ? _GEN_1959 : grid_127; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2264 = 2'h2 == currentTask ? _GEN_1960 : grid_128; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2265 = 2'h2 == currentTask ? _GEN_1961 : grid_129; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2266 = 2'h2 == currentTask ? _GEN_1962 : grid_130; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2267 = 2'h2 == currentTask ? _GEN_1963 : grid_131; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2268 = 2'h2 == currentTask ? _GEN_1964 : grid_132; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2269 = 2'h2 == currentTask ? _GEN_1965 : grid_133; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2270 = 2'h2 == currentTask ? _GEN_1966 : grid_134; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2271 = 2'h2 == currentTask ? _GEN_1967 : grid_135; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2272 = 2'h2 == currentTask ? _GEN_1968 : grid_136; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2273 = 2'h2 == currentTask ? _GEN_1969 : grid_137; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2274 = 2'h2 == currentTask ? _GEN_1970 : grid_138; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2275 = 2'h2 == currentTask ? _GEN_1971 : grid_139; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2276 = 2'h2 == currentTask ? _GEN_1972 : grid_140; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2277 = 2'h2 == currentTask ? _GEN_1973 : grid_141; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2278 = 2'h2 == currentTask ? _GEN_1974 : grid_142; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2279 = 2'h2 == currentTask ? _GEN_1975 : grid_143; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2280 = 2'h2 == currentTask ? _GEN_1976 : grid_144; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2281 = 2'h2 == currentTask ? _GEN_1977 : grid_145; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2282 = 2'h2 == currentTask ? _GEN_1978 : grid_146; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2283 = 2'h2 == currentTask ? _GEN_1979 : grid_147; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2284 = 2'h2 == currentTask ? _GEN_1980 : grid_148; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2285 = 2'h2 == currentTask ? _GEN_1981 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2286 = 2'h2 == currentTask ? _GEN_1982 : grid_150; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2287 = 2'h2 == currentTask ? _GEN_1983 : grid_151; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2288 = 2'h2 == currentTask ? _GEN_1984 : grid_152; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2289 = 2'h2 == currentTask ? _GEN_1985 : grid_153; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2290 = 2'h2 == currentTask ? _GEN_1986 : grid_154; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2291 = 2'h2 == currentTask ? _GEN_1987 : grid_155; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2292 = 2'h2 == currentTask ? _GEN_1988 : grid_156; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2293 = 2'h2 == currentTask ? _GEN_1989 : grid_157; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2294 = 2'h2 == currentTask ? _GEN_1990 : grid_158; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2295 = 2'h2 == currentTask ? _GEN_1991 : grid_159; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2296 = 2'h2 == currentTask ? _GEN_1992 : grid_160; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2297 = 2'h2 == currentTask ? _GEN_1993 : grid_161; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2298 = 2'h2 == currentTask ? _GEN_1994 : grid_162; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2299 = 2'h2 == currentTask ? _GEN_1995 : grid_163; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2300 = 2'h2 == currentTask ? _GEN_1996 : grid_164; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2301 = 2'h2 == currentTask ? _GEN_1997 : grid_165; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2302 = 2'h2 == currentTask ? _GEN_1998 : grid_166; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2303 = 2'h2 == currentTask ? _GEN_1999 : grid_167; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2304 = 2'h2 == currentTask ? _GEN_2000 : grid_168; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2305 = 2'h2 == currentTask ? _GEN_2001 : grid_169; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2306 = 2'h2 == currentTask ? _GEN_2002 : grid_170; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2307 = 2'h2 == currentTask ? _GEN_2003 : grid_171; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2308 = 2'h2 == currentTask ? _GEN_2004 : grid_172; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2309 = 2'h2 == currentTask ? _GEN_2005 : grid_173; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2310 = 2'h2 == currentTask ? _GEN_2006 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2311 = 2'h2 == currentTask ? _GEN_2007 : grid_175; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2312 = 2'h2 == currentTask ? _GEN_2008 : grid_176; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2313 = 2'h2 == currentTask ? _GEN_2009 : grid_177; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2314 = 2'h2 == currentTask ? _GEN_2010 : grid_178; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2315 = 2'h2 == currentTask ? _GEN_2011 : grid_179; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2316 = 2'h2 == currentTask ? _GEN_2012 : grid_180; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2317 = 2'h2 == currentTask ? _GEN_2013 : grid_181; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2318 = 2'h2 == currentTask ? _GEN_2014 : grid_182; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2319 = 2'h2 == currentTask ? _GEN_2015 : grid_183; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2320 = 2'h2 == currentTask ? _GEN_2016 : grid_184; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2321 = 2'h2 == currentTask ? _GEN_2017 : grid_185; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2322 = 2'h2 == currentTask ? _GEN_2018 : grid_186; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2323 = 2'h2 == currentTask ? _GEN_2019 : grid_187; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2324 = 2'h2 == currentTask ? _GEN_2020 : grid_188; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2325 = 2'h2 == currentTask ? _GEN_2021 : grid_189; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2326 = 2'h2 == currentTask ? _GEN_2022 : grid_190; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2327 = 2'h2 == currentTask ? _GEN_2023 : grid_191; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2328 = 2'h2 == currentTask ? _GEN_2024 : grid_192; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2329 = 2'h2 == currentTask ? _GEN_2025 : grid_193; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2330 = 2'h2 == currentTask ? _GEN_2026 : grid_194; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2331 = 2'h2 == currentTask ? _GEN_2027 : grid_195; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2332 = 2'h2 == currentTask ? _GEN_2028 : grid_196; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2333 = 2'h2 == currentTask ? _GEN_2029 : grid_197; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2334 = 2'h2 == currentTask ? _GEN_2030 : grid_198; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2335 = 2'h2 == currentTask ? _GEN_2031 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2336 = 2'h2 == currentTask ? _GEN_2032 : grid_200; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2337 = 2'h2 == currentTask ? _GEN_2033 : grid_201; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2338 = 2'h2 == currentTask ? _GEN_2034 : grid_202; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2339 = 2'h2 == currentTask ? _GEN_2035 : grid_203; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2340 = 2'h2 == currentTask ? _GEN_2036 : grid_204; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2341 = 2'h2 == currentTask ? _GEN_2037 : grid_205; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2342 = 2'h2 == currentTask ? _GEN_2038 : grid_206; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2343 = 2'h2 == currentTask ? _GEN_2039 : grid_207; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2344 = 2'h2 == currentTask ? _GEN_2040 : grid_208; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2345 = 2'h2 == currentTask ? _GEN_2041 : grid_209; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2346 = 2'h2 == currentTask ? _GEN_2042 : grid_210; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2347 = 2'h2 == currentTask ? _GEN_2043 : grid_211; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2348 = 2'h2 == currentTask ? _GEN_2044 : grid_212; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2349 = 2'h2 == currentTask ? _GEN_2045 : grid_213; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2350 = 2'h2 == currentTask ? _GEN_2046 : grid_214; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2351 = 2'h2 == currentTask ? _GEN_2047 : grid_215; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2352 = 2'h2 == currentTask ? _GEN_2048 : grid_216; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2353 = 2'h2 == currentTask ? _GEN_2049 : grid_217; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2354 = 2'h2 == currentTask ? _GEN_2050 : grid_218; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2355 = 2'h2 == currentTask ? _GEN_2051 : grid_219; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2356 = 2'h2 == currentTask ? _GEN_2052 : grid_220; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2357 = 2'h2 == currentTask ? _GEN_2053 : grid_221; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2358 = 2'h2 == currentTask ? _GEN_2054 : grid_222; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2359 = 2'h2 == currentTask ? _GEN_2055 : grid_223; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2360 = 2'h2 == currentTask ? _GEN_2056 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2361 = 2'h2 == currentTask ? _GEN_2057 : grid_225; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2362 = 2'h2 == currentTask ? _GEN_2058 : grid_226; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2363 = 2'h2 == currentTask ? _GEN_2059 : grid_227; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2364 = 2'h2 == currentTask ? _GEN_2060 : grid_228; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2365 = 2'h2 == currentTask ? _GEN_2061 : grid_229; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2366 = 2'h2 == currentTask ? _GEN_2062 : grid_230; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2367 = 2'h2 == currentTask ? _GEN_2063 : grid_231; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2368 = 2'h2 == currentTask ? _GEN_2064 : grid_232; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2369 = 2'h2 == currentTask ? _GEN_2065 : grid_233; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2370 = 2'h2 == currentTask ? _GEN_2066 : grid_234; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2371 = 2'h2 == currentTask ? _GEN_2067 : grid_235; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2372 = 2'h2 == currentTask ? _GEN_2068 : grid_236; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2373 = 2'h2 == currentTask ? _GEN_2069 : grid_237; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2374 = 2'h2 == currentTask ? _GEN_2070 : grid_238; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2375 = 2'h2 == currentTask ? _GEN_2071 : grid_239; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2376 = 2'h2 == currentTask ? _GEN_2072 : grid_240; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2377 = 2'h2 == currentTask ? _GEN_2073 : grid_241; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2378 = 2'h2 == currentTask ? _GEN_2074 : grid_242; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2379 = 2'h2 == currentTask ? _GEN_2075 : grid_243; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2380 = 2'h2 == currentTask ? _GEN_2076 : grid_244; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2381 = 2'h2 == currentTask ? _GEN_2077 : grid_245; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2382 = 2'h2 == currentTask ? _GEN_2078 : grid_246; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2383 = 2'h2 == currentTask ? _GEN_2079 : grid_247; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2384 = 2'h2 == currentTask ? _GEN_2080 : grid_248; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2385 = 2'h2 == currentTask ? _GEN_2081 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2386 = 2'h2 == currentTask ? _GEN_2082 : grid_250; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2387 = 2'h2 == currentTask ? _GEN_2083 : grid_251; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2388 = 2'h2 == currentTask ? _GEN_2084 : grid_252; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2389 = 2'h2 == currentTask ? _GEN_2085 : grid_253; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2390 = 2'h2 == currentTask ? _GEN_2086 : grid_254; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2391 = 2'h2 == currentTask ? _GEN_2087 : grid_255; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2392 = 2'h2 == currentTask ? _GEN_2088 : grid_256; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2393 = 2'h2 == currentTask ? _GEN_2089 : grid_257; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2394 = 2'h2 == currentTask ? _GEN_2090 : grid_258; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2395 = 2'h2 == currentTask ? _GEN_2091 : grid_259; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2396 = 2'h2 == currentTask ? _GEN_2092 : grid_260; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2397 = 2'h2 == currentTask ? _GEN_2093 : grid_261; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2398 = 2'h2 == currentTask ? _GEN_2094 : grid_262; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2399 = 2'h2 == currentTask ? _GEN_2095 : grid_263; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2400 = 2'h2 == currentTask ? _GEN_2096 : grid_264; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2401 = 2'h2 == currentTask ? _GEN_2097 : grid_265; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2402 = 2'h2 == currentTask ? _GEN_2098 : grid_266; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2403 = 2'h2 == currentTask ? _GEN_2099 : grid_267; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2404 = 2'h2 == currentTask ? _GEN_2100 : grid_268; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2405 = 2'h2 == currentTask ? _GEN_2101 : grid_269; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2406 = 2'h2 == currentTask ? _GEN_2102 : grid_270; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2407 = 2'h2 == currentTask ? _GEN_2103 : grid_271; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2408 = 2'h2 == currentTask ? _GEN_2104 : grid_272; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2409 = 2'h2 == currentTask ? _GEN_2105 : grid_273; // @[\\src\\main\\scala\\GameLogic.scala 196:27 88:21]
  wire [1:0] _GEN_2410 = 2'h2 == currentTask ? _GEN_2106 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 91:23]
  wire [1:0] _GEN_2411 = 2'h2 == currentTask ? _GEN_2107 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2412 = 2'h2 == currentTask ? _GEN_2108 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2413 = 2'h2 == currentTask ? _GEN_2109 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2414 = 2'h2 == currentTask ? _GEN_2110 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2415 = 2'h2 == currentTask ? _GEN_2111 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2416 = 2'h2 == currentTask ? _GEN_2112 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2417 = 2'h2 == currentTask ? _GEN_2113 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2418 = 2'h2 == currentTask ? _GEN_2114 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2419 = 2'h2 == currentTask ? _GEN_2115 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2420 = 2'h2 == currentTask ? _GEN_2116 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2421 = 2'h2 == currentTask ? _GEN_2117 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2422 = 2'h2 == currentTask ? _GEN_2118 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2423 = 2'h2 == currentTask ? _GEN_2119 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2424 = 2'h2 == currentTask ? _GEN_2120 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2425 = 2'h2 == currentTask ? _GEN_2121 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2426 = 2'h2 == currentTask ? _GEN_2122 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2427 = 2'h2 == currentTask ? _GEN_2123 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2428 = 2'h2 == currentTask ? _GEN_2124 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2429 = 2'h2 == currentTask ? _GEN_2125 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2430 = 2'h2 == currentTask ? _GEN_2126 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2431 = 2'h2 == currentTask ? _GEN_2127 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2432 = 2'h2 == currentTask ? _GEN_2128 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2433 = 2'h2 == currentTask ? _GEN_2129 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2434 = 2'h2 == currentTask ? _GEN_2130 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [1:0] _GEN_2435 = 2'h2 == currentTask ? _GEN_2131 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 196:27 96:21]
  wire [10:0] _GEN_2437 = 2'h1 == currentTask ? $signed(_posToGridIndex_io_xPos_T_2) : $signed(11'sh0); // @[\\src\\main\\scala\\GameLogic.scala 124:26 196:27 199:34]
  wire [9:0] _GEN_2438 = 2'h1 == currentTask ? $signed(_posToGridIndex_io_yPos_T_2) : $signed(10'sh0); // @[\\src\\main\\scala\\GameLogic.scala 125:26 196:27 200:34]
  wire [4:0] _GEN_2741 = 2'h1 == currentTask ? blockLogic_io_tileNumber : _GEN_2135; // @[\\src\\main\\scala\\GameLogic.scala 196:27 204:34]
  wire [10:0] _GEN_2749 = 2'h1 == currentTask ? posToIndex_io_index : {{2'd0}, _GEN_2134}; // @[\\src\\main\\scala\\GameLogic.scala 196:27 216:37]
  wire [2:0] _GEN_2751 = newPiece ? rnd : blockType; // @[\\src\\main\\scala\\GameLogic.scala 249:22 250:19 157:26]
  wire  _GEN_2752 = newPiece ? 1'h0 : newPiece; // @[\\src\\main\\scala\\GameLogic.scala 249:22 251:18 165:25]
  wire [6:0] _moveCnt_T_1 = moveCnt + 7'h1; // @[\\src\\main\\scala\\GameLogic.scala 258:39]
  wire [6:0] _GEN_2753 = moveCnt >= speedThreshold ? 7'h0 : _moveCnt_T_1; // @[\\src\\main\\scala\\GameLogic.scala 254:39 255:17 258:28]
  wire [10:0] fallen = moveCnt >= speedThreshold ? $signed(11'sh1) : $signed(11'sh0); // @[\\src\\main\\scala\\GameLogic.scala 254:39 256:16 245:28]
  wire [9:0] _GEN_2755 = io_btnR ? $signed(-10'sh1) : $signed(10'sh0); // @[\\src\\main\\scala\\GameLogic.scala 262:26 246:27 262:34]
  wire [9:0] moved = io_btnL ? $signed(10'sh1) : $signed(_GEN_2755); // @[\\src\\main\\scala\\GameLogic.scala 261:{21,29}]
  wire [10:0] fallenX = $signed(blockXReg) + $signed(fallen); // @[\\src\\main\\scala\\GameLogic.scala 264:31]
  wire [9:0] movedY = $signed(blockYReg) + $signed(moved); // @[\\src\\main\\scala\\GameLogic.scala 268:30]
  wire  _T_13 = io_btnU & upRelease; // @[\\src\\main\\scala\\GameLogic.scala 280:22]
  wire [1:0] _rotation_T_1 = rotation + 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 284:32]
  wire [1:0] _GEN_2757 = _T_13 ? _rotation_T_1 : rotation; // @[\\src\\main\\scala\\GameLogic.scala 283:43 284:20 147:25]
  wire  _GEN_2758 = _T_13 ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameLogic.scala 283:43 285:21 286:33]
  wire [1:0] _GEN_2759 = io_btnU & upRelease & rotation == 2'h3 ? 2'h0 : _GEN_2757; // @[\\src\\main\\scala\\GameLogic.scala 280:56 281:20]
  wire  _GEN_2760 = io_btnU & upRelease & rotation == 2'h3 ? upRelease : _GEN_2758; // @[\\src\\main\\scala\\GameLogic.scala 149:26 280:56]
  wire [10:0] _GEN_2761 = ~fallDetector_io_isCollision ? $signed(fallenX) : $signed(blockXReg); // @[\\src\\main\\scala\\GameLogic.scala 287:49 288:19 102:26]
  wire [1:0] _GEN_2763 = ~fallDetector_io_isCollision ? 2'h3 : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 243:31 287:49 292:19]
  wire [1:0] _GEN_2764 = ~fallDetector_io_isCollision ? currentTask : 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 287:49 293:21 80:28]
  wire [10:0] _GEN_2765 = ~movementDetector_io_isCollision ? $signed(fallenX) : $signed(_GEN_2761); // @[\\src\\main\\scala\\GameLogic.scala 277:47 278:19]
  wire [9:0] _GEN_2766 = ~movementDetector_io_isCollision ? $signed(movedY) : $signed(blockYReg); // @[\\src\\main\\scala\\GameLogic.scala 277:47 279:19]
  wire [1:0] _GEN_2767 = ~movementDetector_io_isCollision ? _GEN_2759 : rotation; // @[\\src\\main\\scala\\GameLogic.scala 147:25 277:47]
  wire  _GEN_2768 = ~movementDetector_io_isCollision ? _GEN_2760 : upRelease; // @[\\src\\main\\scala\\GameLogic.scala 149:26 277:47]
  wire [1:0] nextState = ~movementDetector_io_isCollision ? 2'h3 : _GEN_2763; // @[\\src\\main\\scala\\GameLogic.scala 243:31 277:47]
  wire [1:0] _GEN_2770 = ~movementDetector_io_isCollision ? currentTask : _GEN_2764; // @[\\src\\main\\scala\\GameLogic.scala 277:47 80:28]
  wire [3:0] _GEN_2771 = io_btnU ? $signed(blockLogic_io_nextOffsetX_0) : $signed(blockLogic_io_activeOffsetX_0); // @[\\src\\main\\scala\\GameLogic.scala 310:21 299:36 311:38]
  wire [3:0] _GEN_2772 = io_btnU ? $signed(blockLogic_io_nextOffsetX_1) : $signed(blockLogic_io_activeOffsetX_1); // @[\\src\\main\\scala\\GameLogic.scala 310:21 299:36 311:38]
  wire [3:0] _GEN_2773 = io_btnU ? $signed(blockLogic_io_nextOffsetX_2) : $signed(blockLogic_io_activeOffsetX_2); // @[\\src\\main\\scala\\GameLogic.scala 310:21 299:36 311:38]
  wire [3:0] _GEN_2774 = io_btnU ? $signed(blockLogic_io_nextOffsetX_3) : $signed(blockLogic_io_activeOffsetX_3); // @[\\src\\main\\scala\\GameLogic.scala 310:21 299:36 311:38]
  wire [3:0] _GEN_2775 = io_btnU ? $signed(blockLogic_io_nextOffsetY_0) : $signed(blockLogic_io_activeOffsetY_0); // @[\\src\\main\\scala\\GameLogic.scala 310:21 300:36 312:38]
  wire [3:0] _GEN_2776 = io_btnU ? $signed(blockLogic_io_nextOffsetY_1) : $signed(blockLogic_io_activeOffsetY_1); // @[\\src\\main\\scala\\GameLogic.scala 310:21 300:36 312:38]
  wire [3:0] _GEN_2777 = io_btnU ? $signed(blockLogic_io_nextOffsetY_2) : $signed(blockLogic_io_activeOffsetY_2); // @[\\src\\main\\scala\\GameLogic.scala 310:21 300:36 312:38]
  wire [3:0] _GEN_2778 = io_btnU ? $signed(blockLogic_io_nextOffsetY_3) : $signed(blockLogic_io_activeOffsetY_3); // @[\\src\\main\\scala\\GameLogic.scala 310:21 300:36 312:38]
  wire [1:0] _GEN_2780 = 2'h3 == stateReg ? 2'h0 : stateReg; // @[\\src\\main\\scala\\GameLogic.scala 186:20 319:16 137:25]
  wire [10:0] _GEN_2785 = 2'h2 == stateReg ? $signed(fallenX) : $signed(blockXReg); // @[\\src\\main\\scala\\GameLogic.scala 186:20 108:24 271:28]
  wire [9:0] _GEN_2788 = 2'h2 == stateReg ? $signed(movedY) : $signed(blockYReg); // @[\\src\\main\\scala\\GameLogic.scala 186:20 115:28 274:32]
  wire  _GEN_2792 = 2'h2 == stateReg ? _GEN_2768 : upRelease; // @[\\src\\main\\scala\\GameLogic.scala 186:20 149:26]
  wire [3:0] _GEN_2794 = 2'h2 == stateReg ? $signed(blockLogic_io_activeOffsetX_0) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28 297:32]
  wire [3:0] _GEN_2795 = 2'h2 == stateReg ? $signed(blockLogic_io_activeOffsetX_1) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28 297:32]
  wire [3:0] _GEN_2796 = 2'h2 == stateReg ? $signed(blockLogic_io_activeOffsetX_2) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28 297:32]
  wire [3:0] _GEN_2797 = 2'h2 == stateReg ? $signed(blockLogic_io_activeOffsetX_3) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28 297:32]
  wire [3:0] _GEN_2798 = 2'h2 == stateReg ? $signed(blockLogic_io_activeOffsetY_0) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28 298:32]
  wire [3:0] _GEN_2799 = 2'h2 == stateReg ? $signed(blockLogic_io_activeOffsetY_1) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28 298:32]
  wire [3:0] _GEN_2800 = 2'h2 == stateReg ? $signed(blockLogic_io_activeOffsetY_2) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28 298:32]
  wire [3:0] _GEN_2801 = 2'h2 == stateReg ? $signed(blockLogic_io_activeOffsetY_3) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28 298:32]
  wire [3:0] _GEN_2802 = 2'h2 == stateReg ? $signed(_GEN_2771) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  wire [3:0] _GEN_2803 = 2'h2 == stateReg ? $signed(_GEN_2772) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  wire [3:0] _GEN_2804 = 2'h2 == stateReg ? $signed(_GEN_2773) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  wire [3:0] _GEN_2805 = 2'h2 == stateReg ? $signed(_GEN_2774) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  wire [3:0] _GEN_2806 = 2'h2 == stateReg ? $signed(_GEN_2775) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  wire [3:0] _GEN_2807 = 2'h2 == stateReg ? $signed(_GEN_2776) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  wire [3:0] _GEN_2808 = 2'h2 == stateReg ? $signed(_GEN_2777) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  wire [3:0] _GEN_2809 = 2'h2 == stateReg ? $signed(_GEN_2778) : $signed(4'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  wire  _GEN_2811 = 2'h2 == stateReg ? 1'h0 : 2'h3 == stateReg; // @[\\src\\main\\scala\\GameLogic.scala 186:20 133:22]
  wire [10:0] _GEN_2813 = 2'h1 == stateReg ? $signed(_GEN_2437) : $signed(11'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 124:26]
  wire [9:0] _GEN_2814 = 2'h1 == stateReg ? $signed(_GEN_2438) : $signed(10'sh0); // @[\\src\\main\\scala\\GameLogic.scala 186:20 125:26]
  wire [4:0] _GEN_3117 = 2'h1 == stateReg ? _GEN_2741 : 5'h0; // @[\\src\\main\\scala\\GameLogic.scala 186:20 128:26]
  wire [10:0] _GEN_3125 = 2'h1 == stateReg ? _GEN_2749 : 11'h0; // @[\\src\\main\\scala\\GameLogic.scala 186:20 129:29]
  wire  _GEN_3127 = 2'h1 == stateReg ? 1'h0 : 2'h2 == stateReg; // @[\\src\\main\\scala\\GameLogic.scala 186:20 76:19]
  wire [10:0] _GEN_3130 = 2'h1 == stateReg ? $signed(blockXReg) : $signed(_GEN_2785); // @[\\src\\main\\scala\\GameLogic.scala 186:20 108:24]
  wire [9:0] _GEN_3133 = 2'h1 == stateReg ? $signed(blockYReg) : $signed(_GEN_2788); // @[\\src\\main\\scala\\GameLogic.scala 186:20 115:28]
  wire  _GEN_3134 = 2'h1 == stateReg ? upRelease : _GEN_2792; // @[\\src\\main\\scala\\GameLogic.scala 186:20 149:26]
  wire [3:0] _GEN_3135 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2794); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28]
  wire [3:0] _GEN_3136 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2795); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28]
  wire [3:0] _GEN_3137 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2796); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28]
  wire [3:0] _GEN_3138 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2797); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28]
  wire [3:0] _GEN_3139 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2798); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28]
  wire [3:0] _GEN_3140 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2799); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28]
  wire [3:0] _GEN_3141 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2800); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28]
  wire [3:0] _GEN_3142 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2801); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28]
  wire [3:0] _GEN_3143 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2802); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  wire [3:0] _GEN_3144 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2803); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  wire [3:0] _GEN_3145 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2804); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  wire [3:0] _GEN_3146 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2805); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  wire [3:0] _GEN_3147 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2806); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  wire [3:0] _GEN_3148 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2807); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  wire [3:0] _GEN_3149 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2808); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  wire [3:0] _GEN_3150 = 2'h1 == stateReg ? $signed(4'sh0) : $signed(_GEN_2809); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  wire  _GEN_3151 = 2'h1 == stateReg ? 1'h0 : _GEN_2811; // @[\\src\\main\\scala\\GameLogic.scala 186:20 133:22]
  wire  _GEN_3474 = 2'h0 == stateReg ? upRelease : _GEN_3134; // @[\\src\\main\\scala\\GameLogic.scala 186:20 149:26]
  CollisionDetector fallDetector ( // @[\\src\\main\\scala\\GameLogic.scala 106:28]
    .io_grid_0(fallDetector_io_grid_0),
    .io_grid_1(fallDetector_io_grid_1),
    .io_grid_2(fallDetector_io_grid_2),
    .io_grid_3(fallDetector_io_grid_3),
    .io_grid_4(fallDetector_io_grid_4),
    .io_grid_5(fallDetector_io_grid_5),
    .io_grid_6(fallDetector_io_grid_6),
    .io_grid_7(fallDetector_io_grid_7),
    .io_grid_8(fallDetector_io_grid_8),
    .io_grid_9(fallDetector_io_grid_9),
    .io_grid_10(fallDetector_io_grid_10),
    .io_grid_11(fallDetector_io_grid_11),
    .io_grid_12(fallDetector_io_grid_12),
    .io_grid_13(fallDetector_io_grid_13),
    .io_grid_14(fallDetector_io_grid_14),
    .io_grid_15(fallDetector_io_grid_15),
    .io_grid_16(fallDetector_io_grid_16),
    .io_grid_17(fallDetector_io_grid_17),
    .io_grid_18(fallDetector_io_grid_18),
    .io_grid_19(fallDetector_io_grid_19),
    .io_grid_20(fallDetector_io_grid_20),
    .io_grid_21(fallDetector_io_grid_21),
    .io_grid_22(fallDetector_io_grid_22),
    .io_grid_23(fallDetector_io_grid_23),
    .io_grid_24(fallDetector_io_grid_24),
    .io_grid_25(fallDetector_io_grid_25),
    .io_grid_26(fallDetector_io_grid_26),
    .io_grid_27(fallDetector_io_grid_27),
    .io_grid_28(fallDetector_io_grid_28),
    .io_grid_29(fallDetector_io_grid_29),
    .io_grid_30(fallDetector_io_grid_30),
    .io_grid_31(fallDetector_io_grid_31),
    .io_grid_32(fallDetector_io_grid_32),
    .io_grid_33(fallDetector_io_grid_33),
    .io_grid_34(fallDetector_io_grid_34),
    .io_grid_35(fallDetector_io_grid_35),
    .io_grid_36(fallDetector_io_grid_36),
    .io_grid_37(fallDetector_io_grid_37),
    .io_grid_38(fallDetector_io_grid_38),
    .io_grid_39(fallDetector_io_grid_39),
    .io_grid_40(fallDetector_io_grid_40),
    .io_grid_41(fallDetector_io_grid_41),
    .io_grid_42(fallDetector_io_grid_42),
    .io_grid_43(fallDetector_io_grid_43),
    .io_grid_44(fallDetector_io_grid_44),
    .io_grid_45(fallDetector_io_grid_45),
    .io_grid_46(fallDetector_io_grid_46),
    .io_grid_47(fallDetector_io_grid_47),
    .io_grid_48(fallDetector_io_grid_48),
    .io_grid_49(fallDetector_io_grid_49),
    .io_grid_50(fallDetector_io_grid_50),
    .io_grid_51(fallDetector_io_grid_51),
    .io_grid_52(fallDetector_io_grid_52),
    .io_grid_53(fallDetector_io_grid_53),
    .io_grid_54(fallDetector_io_grid_54),
    .io_grid_55(fallDetector_io_grid_55),
    .io_grid_56(fallDetector_io_grid_56),
    .io_grid_57(fallDetector_io_grid_57),
    .io_grid_58(fallDetector_io_grid_58),
    .io_grid_59(fallDetector_io_grid_59),
    .io_grid_60(fallDetector_io_grid_60),
    .io_grid_61(fallDetector_io_grid_61),
    .io_grid_62(fallDetector_io_grid_62),
    .io_grid_63(fallDetector_io_grid_63),
    .io_grid_64(fallDetector_io_grid_64),
    .io_grid_65(fallDetector_io_grid_65),
    .io_grid_66(fallDetector_io_grid_66),
    .io_grid_67(fallDetector_io_grid_67),
    .io_grid_68(fallDetector_io_grid_68),
    .io_grid_69(fallDetector_io_grid_69),
    .io_grid_70(fallDetector_io_grid_70),
    .io_grid_71(fallDetector_io_grid_71),
    .io_grid_72(fallDetector_io_grid_72),
    .io_grid_73(fallDetector_io_grid_73),
    .io_grid_74(fallDetector_io_grid_74),
    .io_grid_75(fallDetector_io_grid_75),
    .io_grid_76(fallDetector_io_grid_76),
    .io_grid_77(fallDetector_io_grid_77),
    .io_grid_78(fallDetector_io_grid_78),
    .io_grid_79(fallDetector_io_grid_79),
    .io_grid_80(fallDetector_io_grid_80),
    .io_grid_81(fallDetector_io_grid_81),
    .io_grid_82(fallDetector_io_grid_82),
    .io_grid_83(fallDetector_io_grid_83),
    .io_grid_84(fallDetector_io_grid_84),
    .io_grid_85(fallDetector_io_grid_85),
    .io_grid_86(fallDetector_io_grid_86),
    .io_grid_87(fallDetector_io_grid_87),
    .io_grid_88(fallDetector_io_grid_88),
    .io_grid_89(fallDetector_io_grid_89),
    .io_grid_90(fallDetector_io_grid_90),
    .io_grid_91(fallDetector_io_grid_91),
    .io_grid_92(fallDetector_io_grid_92),
    .io_grid_93(fallDetector_io_grid_93),
    .io_grid_94(fallDetector_io_grid_94),
    .io_grid_95(fallDetector_io_grid_95),
    .io_grid_96(fallDetector_io_grid_96),
    .io_grid_97(fallDetector_io_grid_97),
    .io_grid_98(fallDetector_io_grid_98),
    .io_grid_99(fallDetector_io_grid_99),
    .io_grid_100(fallDetector_io_grid_100),
    .io_grid_101(fallDetector_io_grid_101),
    .io_grid_102(fallDetector_io_grid_102),
    .io_grid_103(fallDetector_io_grid_103),
    .io_grid_104(fallDetector_io_grid_104),
    .io_grid_105(fallDetector_io_grid_105),
    .io_grid_106(fallDetector_io_grid_106),
    .io_grid_107(fallDetector_io_grid_107),
    .io_grid_108(fallDetector_io_grid_108),
    .io_grid_109(fallDetector_io_grid_109),
    .io_grid_110(fallDetector_io_grid_110),
    .io_grid_111(fallDetector_io_grid_111),
    .io_grid_112(fallDetector_io_grid_112),
    .io_grid_113(fallDetector_io_grid_113),
    .io_grid_114(fallDetector_io_grid_114),
    .io_grid_115(fallDetector_io_grid_115),
    .io_grid_116(fallDetector_io_grid_116),
    .io_grid_117(fallDetector_io_grid_117),
    .io_grid_118(fallDetector_io_grid_118),
    .io_grid_119(fallDetector_io_grid_119),
    .io_grid_120(fallDetector_io_grid_120),
    .io_grid_121(fallDetector_io_grid_121),
    .io_grid_122(fallDetector_io_grid_122),
    .io_grid_123(fallDetector_io_grid_123),
    .io_grid_124(fallDetector_io_grid_124),
    .io_grid_125(fallDetector_io_grid_125),
    .io_grid_126(fallDetector_io_grid_126),
    .io_grid_127(fallDetector_io_grid_127),
    .io_grid_128(fallDetector_io_grid_128),
    .io_grid_129(fallDetector_io_grid_129),
    .io_grid_130(fallDetector_io_grid_130),
    .io_grid_131(fallDetector_io_grid_131),
    .io_grid_132(fallDetector_io_grid_132),
    .io_grid_133(fallDetector_io_grid_133),
    .io_grid_134(fallDetector_io_grid_134),
    .io_grid_135(fallDetector_io_grid_135),
    .io_grid_136(fallDetector_io_grid_136),
    .io_grid_137(fallDetector_io_grid_137),
    .io_grid_138(fallDetector_io_grid_138),
    .io_grid_139(fallDetector_io_grid_139),
    .io_grid_140(fallDetector_io_grid_140),
    .io_grid_141(fallDetector_io_grid_141),
    .io_grid_142(fallDetector_io_grid_142),
    .io_grid_143(fallDetector_io_grid_143),
    .io_grid_144(fallDetector_io_grid_144),
    .io_grid_145(fallDetector_io_grid_145),
    .io_grid_146(fallDetector_io_grid_146),
    .io_grid_147(fallDetector_io_grid_147),
    .io_grid_148(fallDetector_io_grid_148),
    .io_grid_149(fallDetector_io_grid_149),
    .io_grid_150(fallDetector_io_grid_150),
    .io_grid_151(fallDetector_io_grid_151),
    .io_grid_152(fallDetector_io_grid_152),
    .io_grid_153(fallDetector_io_grid_153),
    .io_grid_154(fallDetector_io_grid_154),
    .io_grid_155(fallDetector_io_grid_155),
    .io_grid_156(fallDetector_io_grid_156),
    .io_grid_157(fallDetector_io_grid_157),
    .io_grid_158(fallDetector_io_grid_158),
    .io_grid_159(fallDetector_io_grid_159),
    .io_grid_160(fallDetector_io_grid_160),
    .io_grid_161(fallDetector_io_grid_161),
    .io_grid_162(fallDetector_io_grid_162),
    .io_grid_163(fallDetector_io_grid_163),
    .io_grid_164(fallDetector_io_grid_164),
    .io_grid_165(fallDetector_io_grid_165),
    .io_grid_166(fallDetector_io_grid_166),
    .io_grid_167(fallDetector_io_grid_167),
    .io_grid_168(fallDetector_io_grid_168),
    .io_grid_169(fallDetector_io_grid_169),
    .io_grid_170(fallDetector_io_grid_170),
    .io_grid_171(fallDetector_io_grid_171),
    .io_grid_172(fallDetector_io_grid_172),
    .io_grid_173(fallDetector_io_grid_173),
    .io_grid_174(fallDetector_io_grid_174),
    .io_grid_175(fallDetector_io_grid_175),
    .io_grid_176(fallDetector_io_grid_176),
    .io_grid_177(fallDetector_io_grid_177),
    .io_grid_178(fallDetector_io_grid_178),
    .io_grid_179(fallDetector_io_grid_179),
    .io_grid_180(fallDetector_io_grid_180),
    .io_grid_181(fallDetector_io_grid_181),
    .io_grid_182(fallDetector_io_grid_182),
    .io_grid_183(fallDetector_io_grid_183),
    .io_grid_184(fallDetector_io_grid_184),
    .io_grid_185(fallDetector_io_grid_185),
    .io_grid_186(fallDetector_io_grid_186),
    .io_grid_187(fallDetector_io_grid_187),
    .io_grid_188(fallDetector_io_grid_188),
    .io_grid_189(fallDetector_io_grid_189),
    .io_grid_190(fallDetector_io_grid_190),
    .io_grid_191(fallDetector_io_grid_191),
    .io_grid_192(fallDetector_io_grid_192),
    .io_grid_193(fallDetector_io_grid_193),
    .io_grid_194(fallDetector_io_grid_194),
    .io_grid_195(fallDetector_io_grid_195),
    .io_grid_196(fallDetector_io_grid_196),
    .io_grid_197(fallDetector_io_grid_197),
    .io_grid_198(fallDetector_io_grid_198),
    .io_grid_199(fallDetector_io_grid_199),
    .io_grid_200(fallDetector_io_grid_200),
    .io_grid_201(fallDetector_io_grid_201),
    .io_grid_202(fallDetector_io_grid_202),
    .io_grid_203(fallDetector_io_grid_203),
    .io_grid_204(fallDetector_io_grid_204),
    .io_grid_205(fallDetector_io_grid_205),
    .io_grid_206(fallDetector_io_grid_206),
    .io_grid_207(fallDetector_io_grid_207),
    .io_grid_208(fallDetector_io_grid_208),
    .io_grid_209(fallDetector_io_grid_209),
    .io_grid_210(fallDetector_io_grid_210),
    .io_grid_211(fallDetector_io_grid_211),
    .io_grid_212(fallDetector_io_grid_212),
    .io_grid_213(fallDetector_io_grid_213),
    .io_grid_214(fallDetector_io_grid_214),
    .io_grid_215(fallDetector_io_grid_215),
    .io_grid_216(fallDetector_io_grid_216),
    .io_grid_217(fallDetector_io_grid_217),
    .io_grid_218(fallDetector_io_grid_218),
    .io_grid_219(fallDetector_io_grid_219),
    .io_grid_220(fallDetector_io_grid_220),
    .io_grid_221(fallDetector_io_grid_221),
    .io_grid_222(fallDetector_io_grid_222),
    .io_grid_223(fallDetector_io_grid_223),
    .io_grid_224(fallDetector_io_grid_224),
    .io_grid_225(fallDetector_io_grid_225),
    .io_grid_226(fallDetector_io_grid_226),
    .io_grid_227(fallDetector_io_grid_227),
    .io_grid_228(fallDetector_io_grid_228),
    .io_grid_229(fallDetector_io_grid_229),
    .io_grid_230(fallDetector_io_grid_230),
    .io_grid_231(fallDetector_io_grid_231),
    .io_grid_232(fallDetector_io_grid_232),
    .io_grid_233(fallDetector_io_grid_233),
    .io_grid_234(fallDetector_io_grid_234),
    .io_grid_235(fallDetector_io_grid_235),
    .io_grid_236(fallDetector_io_grid_236),
    .io_grid_237(fallDetector_io_grid_237),
    .io_grid_238(fallDetector_io_grid_238),
    .io_grid_239(fallDetector_io_grid_239),
    .io_grid_240(fallDetector_io_grid_240),
    .io_grid_241(fallDetector_io_grid_241),
    .io_grid_242(fallDetector_io_grid_242),
    .io_grid_243(fallDetector_io_grid_243),
    .io_grid_244(fallDetector_io_grid_244),
    .io_grid_245(fallDetector_io_grid_245),
    .io_grid_246(fallDetector_io_grid_246),
    .io_grid_247(fallDetector_io_grid_247),
    .io_grid_248(fallDetector_io_grid_248),
    .io_grid_249(fallDetector_io_grid_249),
    .io_grid_250(fallDetector_io_grid_250),
    .io_grid_251(fallDetector_io_grid_251),
    .io_grid_252(fallDetector_io_grid_252),
    .io_grid_253(fallDetector_io_grid_253),
    .io_grid_254(fallDetector_io_grid_254),
    .io_grid_255(fallDetector_io_grid_255),
    .io_grid_256(fallDetector_io_grid_256),
    .io_grid_257(fallDetector_io_grid_257),
    .io_grid_258(fallDetector_io_grid_258),
    .io_grid_259(fallDetector_io_grid_259),
    .io_grid_260(fallDetector_io_grid_260),
    .io_grid_261(fallDetector_io_grid_261),
    .io_grid_262(fallDetector_io_grid_262),
    .io_grid_263(fallDetector_io_grid_263),
    .io_grid_264(fallDetector_io_grid_264),
    .io_grid_265(fallDetector_io_grid_265),
    .io_grid_266(fallDetector_io_grid_266),
    .io_grid_267(fallDetector_io_grid_267),
    .io_grid_268(fallDetector_io_grid_268),
    .io_grid_269(fallDetector_io_grid_269),
    .io_grid_270(fallDetector_io_grid_270),
    .io_grid_271(fallDetector_io_grid_271),
    .io_grid_272(fallDetector_io_grid_272),
    .io_grid_273(fallDetector_io_grid_273),
    .io_grid_274(fallDetector_io_grid_274),
    .io_grid_275(fallDetector_io_grid_275),
    .io_grid_276(fallDetector_io_grid_276),
    .io_grid_277(fallDetector_io_grid_277),
    .io_grid_278(fallDetector_io_grid_278),
    .io_grid_279(fallDetector_io_grid_279),
    .io_grid_280(fallDetector_io_grid_280),
    .io_grid_281(fallDetector_io_grid_281),
    .io_grid_282(fallDetector_io_grid_282),
    .io_grid_283(fallDetector_io_grid_283),
    .io_grid_284(fallDetector_io_grid_284),
    .io_grid_285(fallDetector_io_grid_285),
    .io_grid_286(fallDetector_io_grid_286),
    .io_grid_287(fallDetector_io_grid_287),
    .io_grid_288(fallDetector_io_grid_288),
    .io_grid_289(fallDetector_io_grid_289),
    .io_grid_290(fallDetector_io_grid_290),
    .io_grid_291(fallDetector_io_grid_291),
    .io_grid_292(fallDetector_io_grid_292),
    .io_grid_293(fallDetector_io_grid_293),
    .io_grid_294(fallDetector_io_grid_294),
    .io_grid_295(fallDetector_io_grid_295),
    .io_grid_296(fallDetector_io_grid_296),
    .io_grid_297(fallDetector_io_grid_297),
    .io_grid_298(fallDetector_io_grid_298),
    .io_grid_299(fallDetector_io_grid_299),
    .io_xPos(fallDetector_io_xPos),
    .io_yPos(fallDetector_io_yPos),
    .io_xOffsets_0(fallDetector_io_xOffsets_0),
    .io_xOffsets_1(fallDetector_io_xOffsets_1),
    .io_xOffsets_2(fallDetector_io_xOffsets_2),
    .io_xOffsets_3(fallDetector_io_xOffsets_3),
    .io_yOffsets_0(fallDetector_io_yOffsets_0),
    .io_yOffsets_1(fallDetector_io_yOffsets_1),
    .io_yOffsets_2(fallDetector_io_yOffsets_2),
    .io_yOffsets_3(fallDetector_io_yOffsets_3),
    .io_isCollision(fallDetector_io_isCollision)
  );
  CollisionDetector movementDetector ( // @[\\src\\main\\scala\\GameLogic.scala 112:32]
    .io_grid_0(movementDetector_io_grid_0),
    .io_grid_1(movementDetector_io_grid_1),
    .io_grid_2(movementDetector_io_grid_2),
    .io_grid_3(movementDetector_io_grid_3),
    .io_grid_4(movementDetector_io_grid_4),
    .io_grid_5(movementDetector_io_grid_5),
    .io_grid_6(movementDetector_io_grid_6),
    .io_grid_7(movementDetector_io_grid_7),
    .io_grid_8(movementDetector_io_grid_8),
    .io_grid_9(movementDetector_io_grid_9),
    .io_grid_10(movementDetector_io_grid_10),
    .io_grid_11(movementDetector_io_grid_11),
    .io_grid_12(movementDetector_io_grid_12),
    .io_grid_13(movementDetector_io_grid_13),
    .io_grid_14(movementDetector_io_grid_14),
    .io_grid_15(movementDetector_io_grid_15),
    .io_grid_16(movementDetector_io_grid_16),
    .io_grid_17(movementDetector_io_grid_17),
    .io_grid_18(movementDetector_io_grid_18),
    .io_grid_19(movementDetector_io_grid_19),
    .io_grid_20(movementDetector_io_grid_20),
    .io_grid_21(movementDetector_io_grid_21),
    .io_grid_22(movementDetector_io_grid_22),
    .io_grid_23(movementDetector_io_grid_23),
    .io_grid_24(movementDetector_io_grid_24),
    .io_grid_25(movementDetector_io_grid_25),
    .io_grid_26(movementDetector_io_grid_26),
    .io_grid_27(movementDetector_io_grid_27),
    .io_grid_28(movementDetector_io_grid_28),
    .io_grid_29(movementDetector_io_grid_29),
    .io_grid_30(movementDetector_io_grid_30),
    .io_grid_31(movementDetector_io_grid_31),
    .io_grid_32(movementDetector_io_grid_32),
    .io_grid_33(movementDetector_io_grid_33),
    .io_grid_34(movementDetector_io_grid_34),
    .io_grid_35(movementDetector_io_grid_35),
    .io_grid_36(movementDetector_io_grid_36),
    .io_grid_37(movementDetector_io_grid_37),
    .io_grid_38(movementDetector_io_grid_38),
    .io_grid_39(movementDetector_io_grid_39),
    .io_grid_40(movementDetector_io_grid_40),
    .io_grid_41(movementDetector_io_grid_41),
    .io_grid_42(movementDetector_io_grid_42),
    .io_grid_43(movementDetector_io_grid_43),
    .io_grid_44(movementDetector_io_grid_44),
    .io_grid_45(movementDetector_io_grid_45),
    .io_grid_46(movementDetector_io_grid_46),
    .io_grid_47(movementDetector_io_grid_47),
    .io_grid_48(movementDetector_io_grid_48),
    .io_grid_49(movementDetector_io_grid_49),
    .io_grid_50(movementDetector_io_grid_50),
    .io_grid_51(movementDetector_io_grid_51),
    .io_grid_52(movementDetector_io_grid_52),
    .io_grid_53(movementDetector_io_grid_53),
    .io_grid_54(movementDetector_io_grid_54),
    .io_grid_55(movementDetector_io_grid_55),
    .io_grid_56(movementDetector_io_grid_56),
    .io_grid_57(movementDetector_io_grid_57),
    .io_grid_58(movementDetector_io_grid_58),
    .io_grid_59(movementDetector_io_grid_59),
    .io_grid_60(movementDetector_io_grid_60),
    .io_grid_61(movementDetector_io_grid_61),
    .io_grid_62(movementDetector_io_grid_62),
    .io_grid_63(movementDetector_io_grid_63),
    .io_grid_64(movementDetector_io_grid_64),
    .io_grid_65(movementDetector_io_grid_65),
    .io_grid_66(movementDetector_io_grid_66),
    .io_grid_67(movementDetector_io_grid_67),
    .io_grid_68(movementDetector_io_grid_68),
    .io_grid_69(movementDetector_io_grid_69),
    .io_grid_70(movementDetector_io_grid_70),
    .io_grid_71(movementDetector_io_grid_71),
    .io_grid_72(movementDetector_io_grid_72),
    .io_grid_73(movementDetector_io_grid_73),
    .io_grid_74(movementDetector_io_grid_74),
    .io_grid_75(movementDetector_io_grid_75),
    .io_grid_76(movementDetector_io_grid_76),
    .io_grid_77(movementDetector_io_grid_77),
    .io_grid_78(movementDetector_io_grid_78),
    .io_grid_79(movementDetector_io_grid_79),
    .io_grid_80(movementDetector_io_grid_80),
    .io_grid_81(movementDetector_io_grid_81),
    .io_grid_82(movementDetector_io_grid_82),
    .io_grid_83(movementDetector_io_grid_83),
    .io_grid_84(movementDetector_io_grid_84),
    .io_grid_85(movementDetector_io_grid_85),
    .io_grid_86(movementDetector_io_grid_86),
    .io_grid_87(movementDetector_io_grid_87),
    .io_grid_88(movementDetector_io_grid_88),
    .io_grid_89(movementDetector_io_grid_89),
    .io_grid_90(movementDetector_io_grid_90),
    .io_grid_91(movementDetector_io_grid_91),
    .io_grid_92(movementDetector_io_grid_92),
    .io_grid_93(movementDetector_io_grid_93),
    .io_grid_94(movementDetector_io_grid_94),
    .io_grid_95(movementDetector_io_grid_95),
    .io_grid_96(movementDetector_io_grid_96),
    .io_grid_97(movementDetector_io_grid_97),
    .io_grid_98(movementDetector_io_grid_98),
    .io_grid_99(movementDetector_io_grid_99),
    .io_grid_100(movementDetector_io_grid_100),
    .io_grid_101(movementDetector_io_grid_101),
    .io_grid_102(movementDetector_io_grid_102),
    .io_grid_103(movementDetector_io_grid_103),
    .io_grid_104(movementDetector_io_grid_104),
    .io_grid_105(movementDetector_io_grid_105),
    .io_grid_106(movementDetector_io_grid_106),
    .io_grid_107(movementDetector_io_grid_107),
    .io_grid_108(movementDetector_io_grid_108),
    .io_grid_109(movementDetector_io_grid_109),
    .io_grid_110(movementDetector_io_grid_110),
    .io_grid_111(movementDetector_io_grid_111),
    .io_grid_112(movementDetector_io_grid_112),
    .io_grid_113(movementDetector_io_grid_113),
    .io_grid_114(movementDetector_io_grid_114),
    .io_grid_115(movementDetector_io_grid_115),
    .io_grid_116(movementDetector_io_grid_116),
    .io_grid_117(movementDetector_io_grid_117),
    .io_grid_118(movementDetector_io_grid_118),
    .io_grid_119(movementDetector_io_grid_119),
    .io_grid_120(movementDetector_io_grid_120),
    .io_grid_121(movementDetector_io_grid_121),
    .io_grid_122(movementDetector_io_grid_122),
    .io_grid_123(movementDetector_io_grid_123),
    .io_grid_124(movementDetector_io_grid_124),
    .io_grid_125(movementDetector_io_grid_125),
    .io_grid_126(movementDetector_io_grid_126),
    .io_grid_127(movementDetector_io_grid_127),
    .io_grid_128(movementDetector_io_grid_128),
    .io_grid_129(movementDetector_io_grid_129),
    .io_grid_130(movementDetector_io_grid_130),
    .io_grid_131(movementDetector_io_grid_131),
    .io_grid_132(movementDetector_io_grid_132),
    .io_grid_133(movementDetector_io_grid_133),
    .io_grid_134(movementDetector_io_grid_134),
    .io_grid_135(movementDetector_io_grid_135),
    .io_grid_136(movementDetector_io_grid_136),
    .io_grid_137(movementDetector_io_grid_137),
    .io_grid_138(movementDetector_io_grid_138),
    .io_grid_139(movementDetector_io_grid_139),
    .io_grid_140(movementDetector_io_grid_140),
    .io_grid_141(movementDetector_io_grid_141),
    .io_grid_142(movementDetector_io_grid_142),
    .io_grid_143(movementDetector_io_grid_143),
    .io_grid_144(movementDetector_io_grid_144),
    .io_grid_145(movementDetector_io_grid_145),
    .io_grid_146(movementDetector_io_grid_146),
    .io_grid_147(movementDetector_io_grid_147),
    .io_grid_148(movementDetector_io_grid_148),
    .io_grid_149(movementDetector_io_grid_149),
    .io_grid_150(movementDetector_io_grid_150),
    .io_grid_151(movementDetector_io_grid_151),
    .io_grid_152(movementDetector_io_grid_152),
    .io_grid_153(movementDetector_io_grid_153),
    .io_grid_154(movementDetector_io_grid_154),
    .io_grid_155(movementDetector_io_grid_155),
    .io_grid_156(movementDetector_io_grid_156),
    .io_grid_157(movementDetector_io_grid_157),
    .io_grid_158(movementDetector_io_grid_158),
    .io_grid_159(movementDetector_io_grid_159),
    .io_grid_160(movementDetector_io_grid_160),
    .io_grid_161(movementDetector_io_grid_161),
    .io_grid_162(movementDetector_io_grid_162),
    .io_grid_163(movementDetector_io_grid_163),
    .io_grid_164(movementDetector_io_grid_164),
    .io_grid_165(movementDetector_io_grid_165),
    .io_grid_166(movementDetector_io_grid_166),
    .io_grid_167(movementDetector_io_grid_167),
    .io_grid_168(movementDetector_io_grid_168),
    .io_grid_169(movementDetector_io_grid_169),
    .io_grid_170(movementDetector_io_grid_170),
    .io_grid_171(movementDetector_io_grid_171),
    .io_grid_172(movementDetector_io_grid_172),
    .io_grid_173(movementDetector_io_grid_173),
    .io_grid_174(movementDetector_io_grid_174),
    .io_grid_175(movementDetector_io_grid_175),
    .io_grid_176(movementDetector_io_grid_176),
    .io_grid_177(movementDetector_io_grid_177),
    .io_grid_178(movementDetector_io_grid_178),
    .io_grid_179(movementDetector_io_grid_179),
    .io_grid_180(movementDetector_io_grid_180),
    .io_grid_181(movementDetector_io_grid_181),
    .io_grid_182(movementDetector_io_grid_182),
    .io_grid_183(movementDetector_io_grid_183),
    .io_grid_184(movementDetector_io_grid_184),
    .io_grid_185(movementDetector_io_grid_185),
    .io_grid_186(movementDetector_io_grid_186),
    .io_grid_187(movementDetector_io_grid_187),
    .io_grid_188(movementDetector_io_grid_188),
    .io_grid_189(movementDetector_io_grid_189),
    .io_grid_190(movementDetector_io_grid_190),
    .io_grid_191(movementDetector_io_grid_191),
    .io_grid_192(movementDetector_io_grid_192),
    .io_grid_193(movementDetector_io_grid_193),
    .io_grid_194(movementDetector_io_grid_194),
    .io_grid_195(movementDetector_io_grid_195),
    .io_grid_196(movementDetector_io_grid_196),
    .io_grid_197(movementDetector_io_grid_197),
    .io_grid_198(movementDetector_io_grid_198),
    .io_grid_199(movementDetector_io_grid_199),
    .io_grid_200(movementDetector_io_grid_200),
    .io_grid_201(movementDetector_io_grid_201),
    .io_grid_202(movementDetector_io_grid_202),
    .io_grid_203(movementDetector_io_grid_203),
    .io_grid_204(movementDetector_io_grid_204),
    .io_grid_205(movementDetector_io_grid_205),
    .io_grid_206(movementDetector_io_grid_206),
    .io_grid_207(movementDetector_io_grid_207),
    .io_grid_208(movementDetector_io_grid_208),
    .io_grid_209(movementDetector_io_grid_209),
    .io_grid_210(movementDetector_io_grid_210),
    .io_grid_211(movementDetector_io_grid_211),
    .io_grid_212(movementDetector_io_grid_212),
    .io_grid_213(movementDetector_io_grid_213),
    .io_grid_214(movementDetector_io_grid_214),
    .io_grid_215(movementDetector_io_grid_215),
    .io_grid_216(movementDetector_io_grid_216),
    .io_grid_217(movementDetector_io_grid_217),
    .io_grid_218(movementDetector_io_grid_218),
    .io_grid_219(movementDetector_io_grid_219),
    .io_grid_220(movementDetector_io_grid_220),
    .io_grid_221(movementDetector_io_grid_221),
    .io_grid_222(movementDetector_io_grid_222),
    .io_grid_223(movementDetector_io_grid_223),
    .io_grid_224(movementDetector_io_grid_224),
    .io_grid_225(movementDetector_io_grid_225),
    .io_grid_226(movementDetector_io_grid_226),
    .io_grid_227(movementDetector_io_grid_227),
    .io_grid_228(movementDetector_io_grid_228),
    .io_grid_229(movementDetector_io_grid_229),
    .io_grid_230(movementDetector_io_grid_230),
    .io_grid_231(movementDetector_io_grid_231),
    .io_grid_232(movementDetector_io_grid_232),
    .io_grid_233(movementDetector_io_grid_233),
    .io_grid_234(movementDetector_io_grid_234),
    .io_grid_235(movementDetector_io_grid_235),
    .io_grid_236(movementDetector_io_grid_236),
    .io_grid_237(movementDetector_io_grid_237),
    .io_grid_238(movementDetector_io_grid_238),
    .io_grid_239(movementDetector_io_grid_239),
    .io_grid_240(movementDetector_io_grid_240),
    .io_grid_241(movementDetector_io_grid_241),
    .io_grid_242(movementDetector_io_grid_242),
    .io_grid_243(movementDetector_io_grid_243),
    .io_grid_244(movementDetector_io_grid_244),
    .io_grid_245(movementDetector_io_grid_245),
    .io_grid_246(movementDetector_io_grid_246),
    .io_grid_247(movementDetector_io_grid_247),
    .io_grid_248(movementDetector_io_grid_248),
    .io_grid_249(movementDetector_io_grid_249),
    .io_grid_250(movementDetector_io_grid_250),
    .io_grid_251(movementDetector_io_grid_251),
    .io_grid_252(movementDetector_io_grid_252),
    .io_grid_253(movementDetector_io_grid_253),
    .io_grid_254(movementDetector_io_grid_254),
    .io_grid_255(movementDetector_io_grid_255),
    .io_grid_256(movementDetector_io_grid_256),
    .io_grid_257(movementDetector_io_grid_257),
    .io_grid_258(movementDetector_io_grid_258),
    .io_grid_259(movementDetector_io_grid_259),
    .io_grid_260(movementDetector_io_grid_260),
    .io_grid_261(movementDetector_io_grid_261),
    .io_grid_262(movementDetector_io_grid_262),
    .io_grid_263(movementDetector_io_grid_263),
    .io_grid_264(movementDetector_io_grid_264),
    .io_grid_265(movementDetector_io_grid_265),
    .io_grid_266(movementDetector_io_grid_266),
    .io_grid_267(movementDetector_io_grid_267),
    .io_grid_268(movementDetector_io_grid_268),
    .io_grid_269(movementDetector_io_grid_269),
    .io_grid_270(movementDetector_io_grid_270),
    .io_grid_271(movementDetector_io_grid_271),
    .io_grid_272(movementDetector_io_grid_272),
    .io_grid_273(movementDetector_io_grid_273),
    .io_grid_274(movementDetector_io_grid_274),
    .io_grid_275(movementDetector_io_grid_275),
    .io_grid_276(movementDetector_io_grid_276),
    .io_grid_277(movementDetector_io_grid_277),
    .io_grid_278(movementDetector_io_grid_278),
    .io_grid_279(movementDetector_io_grid_279),
    .io_grid_280(movementDetector_io_grid_280),
    .io_grid_281(movementDetector_io_grid_281),
    .io_grid_282(movementDetector_io_grid_282),
    .io_grid_283(movementDetector_io_grid_283),
    .io_grid_284(movementDetector_io_grid_284),
    .io_grid_285(movementDetector_io_grid_285),
    .io_grid_286(movementDetector_io_grid_286),
    .io_grid_287(movementDetector_io_grid_287),
    .io_grid_288(movementDetector_io_grid_288),
    .io_grid_289(movementDetector_io_grid_289),
    .io_grid_290(movementDetector_io_grid_290),
    .io_grid_291(movementDetector_io_grid_291),
    .io_grid_292(movementDetector_io_grid_292),
    .io_grid_293(movementDetector_io_grid_293),
    .io_grid_294(movementDetector_io_grid_294),
    .io_grid_295(movementDetector_io_grid_295),
    .io_grid_296(movementDetector_io_grid_296),
    .io_grid_297(movementDetector_io_grid_297),
    .io_grid_298(movementDetector_io_grid_298),
    .io_grid_299(movementDetector_io_grid_299),
    .io_xPos(movementDetector_io_xPos),
    .io_yPos(movementDetector_io_yPos),
    .io_xOffsets_0(movementDetector_io_xOffsets_0),
    .io_xOffsets_1(movementDetector_io_xOffsets_1),
    .io_xOffsets_2(movementDetector_io_xOffsets_2),
    .io_xOffsets_3(movementDetector_io_xOffsets_3),
    .io_yOffsets_0(movementDetector_io_yOffsets_0),
    .io_yOffsets_1(movementDetector_io_yOffsets_1),
    .io_yOffsets_2(movementDetector_io_yOffsets_2),
    .io_yOffsets_3(movementDetector_io_yOffsets_3),
    .io_isCollision(movementDetector_io_isCollision)
  );
  PosToIndex posToIndex ( // @[\\src\\main\\scala\\GameLogic.scala 120:26]
    .io_xPos(posToIndex_io_xPos),
    .io_yPos(posToIndex_io_yPos),
    .io_index(posToIndex_io_index)
  );
  PosToGridIndex posToGridIndex ( // @[\\src\\main\\scala\\GameLogic.scala 123:30]
    .io_xPos(posToGridIndex_io_xPos),
    .io_yPos(posToGridIndex_io_yPos),
    .io_index(posToGridIndex_io_index)
  );
  GameScreen gameScreen ( // @[\\src\\main\\scala\\GameLogic.scala 151:26]
    .clock(gameScreen_clock),
    .reset(gameScreen_reset),
    .io_sw(gameScreen_io_sw),
    .io_viewBoxX(gameScreen_io_viewBoxX),
    .io_viewBoxY(gameScreen_io_viewBoxY),
    .io_staticScreen(gameScreen_io_staticScreen)
  );
  MaxPeriodFibonacciLFSR blockType_prng ( // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
    .clock(blockType_prng_clock),
    .reset(blockType_prng_reset),
    .io_increment(blockType_prng_io_increment),
    .io_out_0(blockType_prng_io_out_0),
    .io_out_1(blockType_prng_io_out_1),
    .io_out_2(blockType_prng_io_out_2)
  );
  MaxPeriodFibonacciLFSR rnd_prng ( // @[src/main/scala/chisel3/util/random/PRNG.scala 91:22]
    .clock(rnd_prng_clock),
    .reset(rnd_prng_reset),
    .io_increment(rnd_prng_io_increment),
    .io_out_0(rnd_prng_io_out_0),
    .io_out_1(rnd_prng_io_out_1),
    .io_out_2(rnd_prng_io_out_2)
  );
  BlockLogic blockLogic ( // @[\\src\\main\\scala\\GameLogic.scala 167:26]
    .io_rotation(blockLogic_io_rotation),
    .io_xPos(blockLogic_io_xPos),
    .io_yPos(blockLogic_io_yPos),
    .io_sel(blockLogic_io_sel),
    .io_spriteXPosition_0(blockLogic_io_spriteXPosition_0),
    .io_spriteXPosition_1(blockLogic_io_spriteXPosition_1),
    .io_spriteXPosition_2(blockLogic_io_spriteXPosition_2),
    .io_spriteXPosition_3(blockLogic_io_spriteXPosition_3),
    .io_spriteXPosition_4(blockLogic_io_spriteXPosition_4),
    .io_spriteXPosition_5(blockLogic_io_spriteXPosition_5),
    .io_spriteXPosition_6(blockLogic_io_spriteXPosition_6),
    .io_spriteXPosition_7(blockLogic_io_spriteXPosition_7),
    .io_spriteXPosition_8(blockLogic_io_spriteXPosition_8),
    .io_spriteXPosition_9(blockLogic_io_spriteXPosition_9),
    .io_spriteXPosition_10(blockLogic_io_spriteXPosition_10),
    .io_spriteXPosition_11(blockLogic_io_spriteXPosition_11),
    .io_spriteXPosition_12(blockLogic_io_spriteXPosition_12),
    .io_spriteXPosition_13(blockLogic_io_spriteXPosition_13),
    .io_spriteXPosition_14(blockLogic_io_spriteXPosition_14),
    .io_spriteXPosition_15(blockLogic_io_spriteXPosition_15),
    .io_spriteXPosition_16(blockLogic_io_spriteXPosition_16),
    .io_spriteXPosition_17(blockLogic_io_spriteXPosition_17),
    .io_spriteXPosition_18(blockLogic_io_spriteXPosition_18),
    .io_spriteXPosition_19(blockLogic_io_spriteXPosition_19),
    .io_spriteXPosition_20(blockLogic_io_spriteXPosition_20),
    .io_spriteXPosition_21(blockLogic_io_spriteXPosition_21),
    .io_spriteXPosition_22(blockLogic_io_spriteXPosition_22),
    .io_spriteXPosition_23(blockLogic_io_spriteXPosition_23),
    .io_spriteXPosition_24(blockLogic_io_spriteXPosition_24),
    .io_spriteXPosition_25(blockLogic_io_spriteXPosition_25),
    .io_spriteXPosition_26(blockLogic_io_spriteXPosition_26),
    .io_spriteXPosition_27(blockLogic_io_spriteXPosition_27),
    .io_spriteYPosition_0(blockLogic_io_spriteYPosition_0),
    .io_spriteYPosition_1(blockLogic_io_spriteYPosition_1),
    .io_spriteYPosition_2(blockLogic_io_spriteYPosition_2),
    .io_spriteYPosition_3(blockLogic_io_spriteYPosition_3),
    .io_spriteYPosition_4(blockLogic_io_spriteYPosition_4),
    .io_spriteYPosition_5(blockLogic_io_spriteYPosition_5),
    .io_spriteYPosition_6(blockLogic_io_spriteYPosition_6),
    .io_spriteYPosition_7(blockLogic_io_spriteYPosition_7),
    .io_spriteYPosition_8(blockLogic_io_spriteYPosition_8),
    .io_spriteYPosition_9(blockLogic_io_spriteYPosition_9),
    .io_spriteYPosition_10(blockLogic_io_spriteYPosition_10),
    .io_spriteYPosition_11(blockLogic_io_spriteYPosition_11),
    .io_spriteYPosition_12(blockLogic_io_spriteYPosition_12),
    .io_spriteYPosition_13(blockLogic_io_spriteYPosition_13),
    .io_spriteYPosition_14(blockLogic_io_spriteYPosition_14),
    .io_spriteYPosition_15(blockLogic_io_spriteYPosition_15),
    .io_spriteYPosition_16(blockLogic_io_spriteYPosition_16),
    .io_spriteYPosition_17(blockLogic_io_spriteYPosition_17),
    .io_spriteYPosition_18(blockLogic_io_spriteYPosition_18),
    .io_spriteYPosition_19(blockLogic_io_spriteYPosition_19),
    .io_spriteYPosition_20(blockLogic_io_spriteYPosition_20),
    .io_spriteYPosition_21(blockLogic_io_spriteYPosition_21),
    .io_spriteYPosition_22(blockLogic_io_spriteYPosition_22),
    .io_spriteYPosition_23(blockLogic_io_spriteYPosition_23),
    .io_spriteYPosition_24(blockLogic_io_spriteYPosition_24),
    .io_spriteYPosition_25(blockLogic_io_spriteYPosition_25),
    .io_spriteYPosition_26(blockLogic_io_spriteYPosition_26),
    .io_spriteYPosition_27(blockLogic_io_spriteYPosition_27),
    .io_spriteVisible_0(blockLogic_io_spriteVisible_0),
    .io_spriteVisible_1(blockLogic_io_spriteVisible_1),
    .io_spriteVisible_2(blockLogic_io_spriteVisible_2),
    .io_spriteVisible_3(blockLogic_io_spriteVisible_3),
    .io_spriteVisible_4(blockLogic_io_spriteVisible_4),
    .io_spriteVisible_5(blockLogic_io_spriteVisible_5),
    .io_spriteVisible_6(blockLogic_io_spriteVisible_6),
    .io_spriteVisible_7(blockLogic_io_spriteVisible_7),
    .io_spriteVisible_8(blockLogic_io_spriteVisible_8),
    .io_spriteVisible_9(blockLogic_io_spriteVisible_9),
    .io_spriteVisible_10(blockLogic_io_spriteVisible_10),
    .io_spriteVisible_11(blockLogic_io_spriteVisible_11),
    .io_spriteVisible_12(blockLogic_io_spriteVisible_12),
    .io_spriteVisible_13(blockLogic_io_spriteVisible_13),
    .io_spriteVisible_14(blockLogic_io_spriteVisible_14),
    .io_spriteVisible_15(blockLogic_io_spriteVisible_15),
    .io_spriteVisible_16(blockLogic_io_spriteVisible_16),
    .io_spriteVisible_17(blockLogic_io_spriteVisible_17),
    .io_spriteVisible_18(blockLogic_io_spriteVisible_18),
    .io_spriteVisible_19(blockLogic_io_spriteVisible_19),
    .io_spriteVisible_20(blockLogic_io_spriteVisible_20),
    .io_spriteVisible_21(blockLogic_io_spriteVisible_21),
    .io_spriteVisible_22(blockLogic_io_spriteVisible_22),
    .io_spriteVisible_23(blockLogic_io_spriteVisible_23),
    .io_spriteVisible_24(blockLogic_io_spriteVisible_24),
    .io_spriteVisible_25(blockLogic_io_spriteVisible_25),
    .io_spriteVisible_26(blockLogic_io_spriteVisible_26),
    .io_spriteVisible_27(blockLogic_io_spriteVisible_27),
    .io_activeOffsetX_0(blockLogic_io_activeOffsetX_0),
    .io_activeOffsetX_1(blockLogic_io_activeOffsetX_1),
    .io_activeOffsetX_2(blockLogic_io_activeOffsetX_2),
    .io_activeOffsetX_3(blockLogic_io_activeOffsetX_3),
    .io_activeOffsetY_0(blockLogic_io_activeOffsetY_0),
    .io_activeOffsetY_1(blockLogic_io_activeOffsetY_1),
    .io_activeOffsetY_2(blockLogic_io_activeOffsetY_2),
    .io_activeOffsetY_3(blockLogic_io_activeOffsetY_3),
    .io_nextOffsetX_0(blockLogic_io_nextOffsetX_0),
    .io_nextOffsetX_1(blockLogic_io_nextOffsetX_1),
    .io_nextOffsetX_2(blockLogic_io_nextOffsetX_2),
    .io_nextOffsetX_3(blockLogic_io_nextOffsetX_3),
    .io_nextOffsetY_0(blockLogic_io_nextOffsetY_0),
    .io_nextOffsetY_1(blockLogic_io_nextOffsetY_1),
    .io_nextOffsetY_2(blockLogic_io_nextOffsetY_2),
    .io_nextOffsetY_3(blockLogic_io_nextOffsetY_3),
    .io_tileNumber(blockLogic_io_tileNumber)
  );
  assign io_led_0 = grid_46[0]; // @[\\src\\main\\scala\\GameLogic.scala 180:13]
  assign io_led_1 = grid_47[0]; // @[\\src\\main\\scala\\GameLogic.scala 181:13]
  assign io_led_2 = grid_48[0]; // @[\\src\\main\\scala\\GameLogic.scala 182:13]
  assign io_led_3 = grid_73[0]; // @[\\src\\main\\scala\\GameLogic.scala 183:13]
  assign io_spriteXPosition_0 = blockLogic_io_spriteXPosition_0; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_1 = blockLogic_io_spriteXPosition_1; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_2 = blockLogic_io_spriteXPosition_2; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_3 = blockLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_4 = blockLogic_io_spriteXPosition_4; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_5 = blockLogic_io_spriteXPosition_5; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_6 = blockLogic_io_spriteXPosition_6; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_7 = blockLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_8 = blockLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_9 = blockLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_10 = blockLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_11 = blockLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_12 = blockLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_13 = blockLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_14 = blockLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_15 = blockLogic_io_spriteXPosition_15; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_16 = blockLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_17 = blockLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_18 = blockLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_19 = blockLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_20 = blockLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_21 = blockLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_22 = blockLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_23 = blockLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_24 = blockLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_25 = blockLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_26 = blockLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteXPosition_27 = blockLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameLogic.scala 173:22]
  assign io_spriteYPosition_0 = blockLogic_io_spriteYPosition_0; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_1 = blockLogic_io_spriteYPosition_1; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_2 = blockLogic_io_spriteYPosition_2; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_3 = blockLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_4 = blockLogic_io_spriteYPosition_4; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_5 = blockLogic_io_spriteYPosition_5; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_6 = blockLogic_io_spriteYPosition_6; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_7 = blockLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_8 = blockLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_9 = blockLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_10 = blockLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_11 = blockLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_12 = blockLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_13 = blockLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_14 = blockLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_15 = blockLogic_io_spriteYPosition_15; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_16 = blockLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_17 = blockLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_18 = blockLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_19 = blockLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_20 = blockLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_21 = blockLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_22 = blockLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_23 = blockLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_24 = blockLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_25 = blockLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_26 = blockLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteYPosition_27 = blockLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameLogic.scala 174:22]
  assign io_spriteVisible_0 = blockLogic_io_spriteVisible_0; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_1 = blockLogic_io_spriteVisible_1; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_2 = blockLogic_io_spriteVisible_2; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_3 = blockLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_4 = blockLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_5 = blockLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_6 = blockLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_7 = blockLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_8 = blockLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_9 = blockLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_10 = blockLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_11 = blockLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_12 = blockLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_13 = blockLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_14 = blockLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_15 = blockLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_16 = blockLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_17 = blockLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_18 = blockLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_19 = blockLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_20 = blockLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_21 = blockLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_22 = blockLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_23 = blockLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_24 = blockLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_25 = blockLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_26 = blockLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_spriteVisible_27 = blockLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameLogic.scala 172:20]
  assign io_viewBoxX = gameScreen_io_viewBoxX; // @[\\src\\main\\scala\\GameLogic.scala 153:15]
  assign io_viewBoxY = gameScreen_io_viewBoxY; // @[\\src\\main\\scala\\GameLogic.scala 154:15]
  assign io_backBufferWriteData = 2'h0 == stateReg ? 5'h0 : _GEN_3117; // @[\\src\\main\\scala\\GameLogic.scala 186:20 128:26]
  assign io_backBufferWriteAddress = 2'h0 == stateReg ? 11'h0 : _GEN_3125; // @[\\src\\main\\scala\\GameLogic.scala 186:20 129:29]
  assign io_backBufferWriteEnable = 2'h0 == stateReg ? 1'h0 : 2'h1 == stateReg & _T_4; // @[\\src\\main\\scala\\GameLogic.scala 186:20 130:28]
  assign io_frameUpdateDone = 2'h0 == stateReg ? 1'h0 : _GEN_3151; // @[\\src\\main\\scala\\GameLogic.scala 186:20 133:22]
  assign io_startTune_0 = 2'h0 == stateReg ? 1'h0 : _GEN_3127; // @[\\src\\main\\scala\\GameLogic.scala 186:20 193:17]
  assign fallDetector_io_grid_0 = {{1'd0}, grid_0}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_1 = {{1'd0}, grid_1}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_2 = {{1'd0}, grid_2}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_3 = {{1'd0}, grid_3}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_4 = {{1'd0}, grid_4}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_5 = {{1'd0}, grid_5}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_6 = {{1'd0}, grid_6}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_7 = {{1'd0}, grid_7}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_8 = {{1'd0}, grid_8}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_9 = {{1'd0}, grid_9}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_10 = {{1'd0}, grid_10}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_11 = {{1'd0}, grid_11}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_12 = {{1'd0}, grid_12}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_13 = {{1'd0}, grid_13}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_14 = {{1'd0}, grid_14}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_15 = {{1'd0}, grid_15}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_16 = {{1'd0}, grid_16}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_17 = {{1'd0}, grid_17}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_18 = {{1'd0}, grid_18}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_19 = {{1'd0}, grid_19}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_20 = {{1'd0}, grid_20}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_21 = {{1'd0}, grid_21}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_22 = {{1'd0}, grid_22}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_23 = {{1'd0}, grid_23}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_24 = {{1'd0}, grid_24}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_25 = {{1'd0}, grid_25}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_26 = {{1'd0}, grid_26}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_27 = {{1'd0}, grid_27}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_28 = {{1'd0}, grid_28}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_29 = {{1'd0}, grid_29}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_30 = {{1'd0}, grid_30}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_31 = {{1'd0}, grid_31}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_32 = {{1'd0}, grid_32}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_33 = {{1'd0}, grid_33}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_34 = {{1'd0}, grid_34}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_35 = {{1'd0}, grid_35}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_36 = {{1'd0}, grid_36}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_37 = {{1'd0}, grid_37}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_38 = {{1'd0}, grid_38}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_39 = {{1'd0}, grid_39}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_40 = {{1'd0}, grid_40}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_41 = {{1'd0}, grid_41}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_42 = {{1'd0}, grid_42}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_43 = {{1'd0}, grid_43}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_44 = {{1'd0}, grid_44}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_45 = {{1'd0}, grid_45}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_46 = {{1'd0}, grid_46}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_47 = {{1'd0}, grid_47}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_48 = {{1'd0}, grid_48}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_49 = {{1'd0}, grid_49}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_50 = {{1'd0}, grid_50}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_51 = {{1'd0}, grid_51}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_52 = {{1'd0}, grid_52}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_53 = {{1'd0}, grid_53}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_54 = {{1'd0}, grid_54}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_55 = {{1'd0}, grid_55}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_56 = {{1'd0}, grid_56}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_57 = {{1'd0}, grid_57}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_58 = {{1'd0}, grid_58}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_59 = {{1'd0}, grid_59}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_60 = {{1'd0}, grid_60}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_61 = {{1'd0}, grid_61}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_62 = {{1'd0}, grid_62}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_63 = {{1'd0}, grid_63}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_64 = {{1'd0}, grid_64}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_65 = {{1'd0}, grid_65}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_66 = {{1'd0}, grid_66}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_67 = {{1'd0}, grid_67}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_68 = {{1'd0}, grid_68}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_69 = {{1'd0}, grid_69}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_70 = {{1'd0}, grid_70}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_71 = {{1'd0}, grid_71}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_72 = {{1'd0}, grid_72}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_73 = {{1'd0}, grid_73}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_74 = {{1'd0}, grid_74}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_75 = {{1'd0}, grid_75}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_76 = {{1'd0}, grid_76}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_77 = {{1'd0}, grid_77}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_78 = {{1'd0}, grid_78}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_79 = {{1'd0}, grid_79}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_80 = {{1'd0}, grid_80}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_81 = {{1'd0}, grid_81}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_82 = {{1'd0}, grid_82}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_83 = {{1'd0}, grid_83}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_84 = {{1'd0}, grid_84}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_85 = {{1'd0}, grid_85}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_86 = {{1'd0}, grid_86}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_87 = {{1'd0}, grid_87}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_88 = {{1'd0}, grid_88}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_89 = {{1'd0}, grid_89}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_90 = {{1'd0}, grid_90}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_91 = {{1'd0}, grid_91}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_92 = {{1'd0}, grid_92}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_93 = {{1'd0}, grid_93}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_94 = {{1'd0}, grid_94}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_95 = {{1'd0}, grid_95}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_96 = {{1'd0}, grid_96}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_97 = {{1'd0}, grid_97}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_98 = {{1'd0}, grid_98}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_99 = {{1'd0}, grid_99}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_100 = {{1'd0}, grid_100}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_101 = {{1'd0}, grid_101}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_102 = {{1'd0}, grid_102}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_103 = {{1'd0}, grid_103}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_104 = {{1'd0}, grid_104}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_105 = {{1'd0}, grid_105}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_106 = {{1'd0}, grid_106}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_107 = {{1'd0}, grid_107}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_108 = {{1'd0}, grid_108}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_109 = {{1'd0}, grid_109}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_110 = {{1'd0}, grid_110}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_111 = {{1'd0}, grid_111}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_112 = {{1'd0}, grid_112}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_113 = {{1'd0}, grid_113}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_114 = {{1'd0}, grid_114}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_115 = {{1'd0}, grid_115}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_116 = {{1'd0}, grid_116}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_117 = {{1'd0}, grid_117}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_118 = {{1'd0}, grid_118}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_119 = {{1'd0}, grid_119}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_120 = {{1'd0}, grid_120}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_121 = {{1'd0}, grid_121}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_122 = {{1'd0}, grid_122}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_123 = {{1'd0}, grid_123}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_124 = {{1'd0}, grid_124}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_125 = {{1'd0}, grid_125}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_126 = {{1'd0}, grid_126}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_127 = {{1'd0}, grid_127}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_128 = {{1'd0}, grid_128}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_129 = {{1'd0}, grid_129}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_130 = {{1'd0}, grid_130}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_131 = {{1'd0}, grid_131}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_132 = {{1'd0}, grid_132}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_133 = {{1'd0}, grid_133}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_134 = {{1'd0}, grid_134}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_135 = {{1'd0}, grid_135}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_136 = {{1'd0}, grid_136}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_137 = {{1'd0}, grid_137}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_138 = {{1'd0}, grid_138}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_139 = {{1'd0}, grid_139}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_140 = {{1'd0}, grid_140}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_141 = {{1'd0}, grid_141}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_142 = {{1'd0}, grid_142}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_143 = {{1'd0}, grid_143}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_144 = {{1'd0}, grid_144}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_145 = {{1'd0}, grid_145}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_146 = {{1'd0}, grid_146}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_147 = {{1'd0}, grid_147}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_148 = {{1'd0}, grid_148}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_149 = {{1'd0}, grid_149}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_150 = {{1'd0}, grid_150}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_151 = {{1'd0}, grid_151}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_152 = {{1'd0}, grid_152}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_153 = {{1'd0}, grid_153}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_154 = {{1'd0}, grid_154}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_155 = {{1'd0}, grid_155}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_156 = {{1'd0}, grid_156}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_157 = {{1'd0}, grid_157}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_158 = {{1'd0}, grid_158}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_159 = {{1'd0}, grid_159}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_160 = {{1'd0}, grid_160}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_161 = {{1'd0}, grid_161}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_162 = {{1'd0}, grid_162}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_163 = {{1'd0}, grid_163}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_164 = {{1'd0}, grid_164}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_165 = {{1'd0}, grid_165}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_166 = {{1'd0}, grid_166}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_167 = {{1'd0}, grid_167}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_168 = {{1'd0}, grid_168}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_169 = {{1'd0}, grid_169}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_170 = {{1'd0}, grid_170}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_171 = {{1'd0}, grid_171}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_172 = {{1'd0}, grid_172}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_173 = {{1'd0}, grid_173}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_174 = {{1'd0}, grid_174}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_175 = {{1'd0}, grid_175}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_176 = {{1'd0}, grid_176}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_177 = {{1'd0}, grid_177}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_178 = {{1'd0}, grid_178}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_179 = {{1'd0}, grid_179}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_180 = {{1'd0}, grid_180}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_181 = {{1'd0}, grid_181}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_182 = {{1'd0}, grid_182}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_183 = {{1'd0}, grid_183}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_184 = {{1'd0}, grid_184}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_185 = {{1'd0}, grid_185}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_186 = {{1'd0}, grid_186}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_187 = {{1'd0}, grid_187}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_188 = {{1'd0}, grid_188}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_189 = {{1'd0}, grid_189}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_190 = {{1'd0}, grid_190}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_191 = {{1'd0}, grid_191}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_192 = {{1'd0}, grid_192}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_193 = {{1'd0}, grid_193}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_194 = {{1'd0}, grid_194}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_195 = {{1'd0}, grid_195}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_196 = {{1'd0}, grid_196}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_197 = {{1'd0}, grid_197}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_198 = {{1'd0}, grid_198}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_199 = {{1'd0}, grid_199}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_200 = {{1'd0}, grid_200}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_201 = {{1'd0}, grid_201}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_202 = {{1'd0}, grid_202}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_203 = {{1'd0}, grid_203}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_204 = {{1'd0}, grid_204}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_205 = {{1'd0}, grid_205}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_206 = {{1'd0}, grid_206}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_207 = {{1'd0}, grid_207}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_208 = {{1'd0}, grid_208}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_209 = {{1'd0}, grid_209}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_210 = {{1'd0}, grid_210}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_211 = {{1'd0}, grid_211}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_212 = {{1'd0}, grid_212}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_213 = {{1'd0}, grid_213}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_214 = {{1'd0}, grid_214}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_215 = {{1'd0}, grid_215}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_216 = {{1'd0}, grid_216}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_217 = {{1'd0}, grid_217}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_218 = {{1'd0}, grid_218}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_219 = {{1'd0}, grid_219}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_220 = {{1'd0}, grid_220}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_221 = {{1'd0}, grid_221}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_222 = {{1'd0}, grid_222}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_223 = {{1'd0}, grid_223}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_224 = {{1'd0}, grid_224}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_225 = {{1'd0}, grid_225}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_226 = {{1'd0}, grid_226}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_227 = {{1'd0}, grid_227}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_228 = {{1'd0}, grid_228}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_229 = {{1'd0}, grid_229}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_230 = {{1'd0}, grid_230}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_231 = {{1'd0}, grid_231}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_232 = {{1'd0}, grid_232}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_233 = {{1'd0}, grid_233}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_234 = {{1'd0}, grid_234}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_235 = {{1'd0}, grid_235}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_236 = {{1'd0}, grid_236}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_237 = {{1'd0}, grid_237}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_238 = {{1'd0}, grid_238}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_239 = {{1'd0}, grid_239}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_240 = {{1'd0}, grid_240}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_241 = {{1'd0}, grid_241}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_242 = {{1'd0}, grid_242}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_243 = {{1'd0}, grid_243}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_244 = {{1'd0}, grid_244}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_245 = {{1'd0}, grid_245}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_246 = {{1'd0}, grid_246}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_247 = {{1'd0}, grid_247}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_248 = {{1'd0}, grid_248}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_249 = {{1'd0}, grid_249}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_250 = {{1'd0}, grid_250}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_251 = {{1'd0}, grid_251}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_252 = {{1'd0}, grid_252}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_253 = {{1'd0}, grid_253}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_254 = {{1'd0}, grid_254}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_255 = {{1'd0}, grid_255}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_256 = {{1'd0}, grid_256}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_257 = {{1'd0}, grid_257}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_258 = {{1'd0}, grid_258}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_259 = {{1'd0}, grid_259}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_260 = {{1'd0}, grid_260}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_261 = {{1'd0}, grid_261}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_262 = {{1'd0}, grid_262}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_263 = {{1'd0}, grid_263}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_264 = {{1'd0}, grid_264}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_265 = {{1'd0}, grid_265}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_266 = {{1'd0}, grid_266}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_267 = {{1'd0}, grid_267}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_268 = {{1'd0}, grid_268}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_269 = {{1'd0}, grid_269}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_270 = {{1'd0}, grid_270}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_271 = {{1'd0}, grid_271}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_272 = {{1'd0}, grid_272}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_273 = {{1'd0}, grid_273}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_274 = {{1'd0}, grid_274}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_275 = {{1'd0}, grid_275}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_276 = {{1'd0}, grid_276}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_277 = {{1'd0}, grid_277}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_278 = {{1'd0}, grid_278}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_279 = {{1'd0}, grid_279}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_280 = {{1'd0}, grid_280}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_281 = {{1'd0}, grid_281}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_282 = {{1'd0}, grid_282}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_283 = {{1'd0}, grid_283}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_284 = {{1'd0}, grid_284}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_285 = {{1'd0}, grid_285}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_286 = {{1'd0}, grid_286}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_287 = {{1'd0}, grid_287}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_288 = {{1'd0}, grid_288}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_289 = {{1'd0}, grid_289}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_290 = {{1'd0}, grid_290}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_291 = {{1'd0}, grid_291}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_292 = {{1'd0}, grid_292}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_293 = {{1'd0}, grid_293}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_294 = {{1'd0}, grid_294}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_295 = {{1'd0}, grid_295}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_296 = {{1'd0}, grid_296}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_297 = {{1'd0}, grid_297}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_298 = {{1'd0}, grid_298}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_grid_299 = {{1'd0}, grid_299}; // @[\\src\\main\\scala\\GameLogic.scala 107:24]
  assign fallDetector_io_xPos = 2'h0 == stateReg ? $signed(blockXReg) : $signed(_GEN_3130); // @[\\src\\main\\scala\\GameLogic.scala 186:20 108:24]
  assign fallDetector_io_yPos = blockYReg; // @[\\src\\main\\scala\\GameLogic.scala 186:20 109:24]
  assign fallDetector_io_xOffsets_0 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3135); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28]
  assign fallDetector_io_xOffsets_1 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3136); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28]
  assign fallDetector_io_xOffsets_2 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3137); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28]
  assign fallDetector_io_xOffsets_3 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3138); // @[\\src\\main\\scala\\GameLogic.scala 186:20 110:28]
  assign fallDetector_io_yOffsets_0 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3139); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28]
  assign fallDetector_io_yOffsets_1 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3140); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28]
  assign fallDetector_io_yOffsets_2 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3141); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28]
  assign fallDetector_io_yOffsets_3 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3142); // @[\\src\\main\\scala\\GameLogic.scala 186:20 111:28]
  assign movementDetector_io_grid_0 = {{1'd0}, grid_0}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_1 = {{1'd0}, grid_1}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_2 = {{1'd0}, grid_2}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_3 = {{1'd0}, grid_3}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_4 = {{1'd0}, grid_4}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_5 = {{1'd0}, grid_5}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_6 = {{1'd0}, grid_6}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_7 = {{1'd0}, grid_7}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_8 = {{1'd0}, grid_8}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_9 = {{1'd0}, grid_9}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_10 = {{1'd0}, grid_10}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_11 = {{1'd0}, grid_11}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_12 = {{1'd0}, grid_12}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_13 = {{1'd0}, grid_13}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_14 = {{1'd0}, grid_14}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_15 = {{1'd0}, grid_15}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_16 = {{1'd0}, grid_16}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_17 = {{1'd0}, grid_17}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_18 = {{1'd0}, grid_18}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_19 = {{1'd0}, grid_19}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_20 = {{1'd0}, grid_20}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_21 = {{1'd0}, grid_21}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_22 = {{1'd0}, grid_22}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_23 = {{1'd0}, grid_23}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_24 = {{1'd0}, grid_24}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_25 = {{1'd0}, grid_25}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_26 = {{1'd0}, grid_26}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_27 = {{1'd0}, grid_27}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_28 = {{1'd0}, grid_28}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_29 = {{1'd0}, grid_29}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_30 = {{1'd0}, grid_30}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_31 = {{1'd0}, grid_31}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_32 = {{1'd0}, grid_32}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_33 = {{1'd0}, grid_33}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_34 = {{1'd0}, grid_34}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_35 = {{1'd0}, grid_35}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_36 = {{1'd0}, grid_36}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_37 = {{1'd0}, grid_37}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_38 = {{1'd0}, grid_38}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_39 = {{1'd0}, grid_39}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_40 = {{1'd0}, grid_40}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_41 = {{1'd0}, grid_41}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_42 = {{1'd0}, grid_42}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_43 = {{1'd0}, grid_43}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_44 = {{1'd0}, grid_44}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_45 = {{1'd0}, grid_45}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_46 = {{1'd0}, grid_46}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_47 = {{1'd0}, grid_47}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_48 = {{1'd0}, grid_48}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_49 = {{1'd0}, grid_49}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_50 = {{1'd0}, grid_50}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_51 = {{1'd0}, grid_51}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_52 = {{1'd0}, grid_52}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_53 = {{1'd0}, grid_53}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_54 = {{1'd0}, grid_54}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_55 = {{1'd0}, grid_55}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_56 = {{1'd0}, grid_56}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_57 = {{1'd0}, grid_57}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_58 = {{1'd0}, grid_58}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_59 = {{1'd0}, grid_59}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_60 = {{1'd0}, grid_60}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_61 = {{1'd0}, grid_61}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_62 = {{1'd0}, grid_62}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_63 = {{1'd0}, grid_63}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_64 = {{1'd0}, grid_64}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_65 = {{1'd0}, grid_65}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_66 = {{1'd0}, grid_66}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_67 = {{1'd0}, grid_67}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_68 = {{1'd0}, grid_68}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_69 = {{1'd0}, grid_69}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_70 = {{1'd0}, grid_70}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_71 = {{1'd0}, grid_71}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_72 = {{1'd0}, grid_72}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_73 = {{1'd0}, grid_73}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_74 = {{1'd0}, grid_74}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_75 = {{1'd0}, grid_75}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_76 = {{1'd0}, grid_76}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_77 = {{1'd0}, grid_77}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_78 = {{1'd0}, grid_78}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_79 = {{1'd0}, grid_79}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_80 = {{1'd0}, grid_80}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_81 = {{1'd0}, grid_81}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_82 = {{1'd0}, grid_82}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_83 = {{1'd0}, grid_83}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_84 = {{1'd0}, grid_84}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_85 = {{1'd0}, grid_85}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_86 = {{1'd0}, grid_86}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_87 = {{1'd0}, grid_87}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_88 = {{1'd0}, grid_88}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_89 = {{1'd0}, grid_89}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_90 = {{1'd0}, grid_90}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_91 = {{1'd0}, grid_91}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_92 = {{1'd0}, grid_92}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_93 = {{1'd0}, grid_93}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_94 = {{1'd0}, grid_94}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_95 = {{1'd0}, grid_95}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_96 = {{1'd0}, grid_96}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_97 = {{1'd0}, grid_97}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_98 = {{1'd0}, grid_98}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_99 = {{1'd0}, grid_99}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_100 = {{1'd0}, grid_100}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_101 = {{1'd0}, grid_101}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_102 = {{1'd0}, grid_102}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_103 = {{1'd0}, grid_103}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_104 = {{1'd0}, grid_104}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_105 = {{1'd0}, grid_105}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_106 = {{1'd0}, grid_106}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_107 = {{1'd0}, grid_107}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_108 = {{1'd0}, grid_108}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_109 = {{1'd0}, grid_109}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_110 = {{1'd0}, grid_110}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_111 = {{1'd0}, grid_111}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_112 = {{1'd0}, grid_112}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_113 = {{1'd0}, grid_113}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_114 = {{1'd0}, grid_114}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_115 = {{1'd0}, grid_115}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_116 = {{1'd0}, grid_116}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_117 = {{1'd0}, grid_117}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_118 = {{1'd0}, grid_118}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_119 = {{1'd0}, grid_119}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_120 = {{1'd0}, grid_120}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_121 = {{1'd0}, grid_121}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_122 = {{1'd0}, grid_122}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_123 = {{1'd0}, grid_123}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_124 = {{1'd0}, grid_124}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_125 = {{1'd0}, grid_125}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_126 = {{1'd0}, grid_126}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_127 = {{1'd0}, grid_127}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_128 = {{1'd0}, grid_128}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_129 = {{1'd0}, grid_129}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_130 = {{1'd0}, grid_130}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_131 = {{1'd0}, grid_131}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_132 = {{1'd0}, grid_132}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_133 = {{1'd0}, grid_133}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_134 = {{1'd0}, grid_134}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_135 = {{1'd0}, grid_135}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_136 = {{1'd0}, grid_136}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_137 = {{1'd0}, grid_137}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_138 = {{1'd0}, grid_138}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_139 = {{1'd0}, grid_139}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_140 = {{1'd0}, grid_140}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_141 = {{1'd0}, grid_141}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_142 = {{1'd0}, grid_142}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_143 = {{1'd0}, grid_143}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_144 = {{1'd0}, grid_144}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_145 = {{1'd0}, grid_145}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_146 = {{1'd0}, grid_146}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_147 = {{1'd0}, grid_147}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_148 = {{1'd0}, grid_148}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_149 = {{1'd0}, grid_149}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_150 = {{1'd0}, grid_150}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_151 = {{1'd0}, grid_151}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_152 = {{1'd0}, grid_152}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_153 = {{1'd0}, grid_153}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_154 = {{1'd0}, grid_154}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_155 = {{1'd0}, grid_155}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_156 = {{1'd0}, grid_156}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_157 = {{1'd0}, grid_157}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_158 = {{1'd0}, grid_158}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_159 = {{1'd0}, grid_159}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_160 = {{1'd0}, grid_160}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_161 = {{1'd0}, grid_161}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_162 = {{1'd0}, grid_162}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_163 = {{1'd0}, grid_163}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_164 = {{1'd0}, grid_164}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_165 = {{1'd0}, grid_165}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_166 = {{1'd0}, grid_166}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_167 = {{1'd0}, grid_167}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_168 = {{1'd0}, grid_168}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_169 = {{1'd0}, grid_169}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_170 = {{1'd0}, grid_170}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_171 = {{1'd0}, grid_171}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_172 = {{1'd0}, grid_172}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_173 = {{1'd0}, grid_173}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_174 = {{1'd0}, grid_174}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_175 = {{1'd0}, grid_175}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_176 = {{1'd0}, grid_176}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_177 = {{1'd0}, grid_177}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_178 = {{1'd0}, grid_178}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_179 = {{1'd0}, grid_179}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_180 = {{1'd0}, grid_180}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_181 = {{1'd0}, grid_181}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_182 = {{1'd0}, grid_182}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_183 = {{1'd0}, grid_183}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_184 = {{1'd0}, grid_184}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_185 = {{1'd0}, grid_185}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_186 = {{1'd0}, grid_186}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_187 = {{1'd0}, grid_187}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_188 = {{1'd0}, grid_188}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_189 = {{1'd0}, grid_189}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_190 = {{1'd0}, grid_190}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_191 = {{1'd0}, grid_191}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_192 = {{1'd0}, grid_192}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_193 = {{1'd0}, grid_193}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_194 = {{1'd0}, grid_194}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_195 = {{1'd0}, grid_195}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_196 = {{1'd0}, grid_196}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_197 = {{1'd0}, grid_197}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_198 = {{1'd0}, grid_198}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_199 = {{1'd0}, grid_199}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_200 = {{1'd0}, grid_200}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_201 = {{1'd0}, grid_201}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_202 = {{1'd0}, grid_202}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_203 = {{1'd0}, grid_203}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_204 = {{1'd0}, grid_204}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_205 = {{1'd0}, grid_205}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_206 = {{1'd0}, grid_206}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_207 = {{1'd0}, grid_207}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_208 = {{1'd0}, grid_208}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_209 = {{1'd0}, grid_209}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_210 = {{1'd0}, grid_210}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_211 = {{1'd0}, grid_211}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_212 = {{1'd0}, grid_212}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_213 = {{1'd0}, grid_213}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_214 = {{1'd0}, grid_214}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_215 = {{1'd0}, grid_215}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_216 = {{1'd0}, grid_216}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_217 = {{1'd0}, grid_217}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_218 = {{1'd0}, grid_218}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_219 = {{1'd0}, grid_219}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_220 = {{1'd0}, grid_220}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_221 = {{1'd0}, grid_221}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_222 = {{1'd0}, grid_222}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_223 = {{1'd0}, grid_223}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_224 = {{1'd0}, grid_224}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_225 = {{1'd0}, grid_225}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_226 = {{1'd0}, grid_226}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_227 = {{1'd0}, grid_227}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_228 = {{1'd0}, grid_228}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_229 = {{1'd0}, grid_229}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_230 = {{1'd0}, grid_230}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_231 = {{1'd0}, grid_231}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_232 = {{1'd0}, grid_232}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_233 = {{1'd0}, grid_233}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_234 = {{1'd0}, grid_234}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_235 = {{1'd0}, grid_235}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_236 = {{1'd0}, grid_236}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_237 = {{1'd0}, grid_237}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_238 = {{1'd0}, grid_238}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_239 = {{1'd0}, grid_239}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_240 = {{1'd0}, grid_240}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_241 = {{1'd0}, grid_241}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_242 = {{1'd0}, grid_242}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_243 = {{1'd0}, grid_243}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_244 = {{1'd0}, grid_244}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_245 = {{1'd0}, grid_245}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_246 = {{1'd0}, grid_246}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_247 = {{1'd0}, grid_247}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_248 = {{1'd0}, grid_248}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_249 = {{1'd0}, grid_249}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_250 = {{1'd0}, grid_250}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_251 = {{1'd0}, grid_251}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_252 = {{1'd0}, grid_252}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_253 = {{1'd0}, grid_253}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_254 = {{1'd0}, grid_254}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_255 = {{1'd0}, grid_255}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_256 = {{1'd0}, grid_256}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_257 = {{1'd0}, grid_257}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_258 = {{1'd0}, grid_258}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_259 = {{1'd0}, grid_259}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_260 = {{1'd0}, grid_260}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_261 = {{1'd0}, grid_261}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_262 = {{1'd0}, grid_262}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_263 = {{1'd0}, grid_263}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_264 = {{1'd0}, grid_264}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_265 = {{1'd0}, grid_265}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_266 = {{1'd0}, grid_266}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_267 = {{1'd0}, grid_267}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_268 = {{1'd0}, grid_268}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_269 = {{1'd0}, grid_269}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_270 = {{1'd0}, grid_270}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_271 = {{1'd0}, grid_271}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_272 = {{1'd0}, grid_272}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_273 = {{1'd0}, grid_273}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_274 = {{1'd0}, grid_274}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_275 = {{1'd0}, grid_275}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_276 = {{1'd0}, grid_276}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_277 = {{1'd0}, grid_277}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_278 = {{1'd0}, grid_278}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_279 = {{1'd0}, grid_279}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_280 = {{1'd0}, grid_280}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_281 = {{1'd0}, grid_281}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_282 = {{1'd0}, grid_282}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_283 = {{1'd0}, grid_283}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_284 = {{1'd0}, grid_284}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_285 = {{1'd0}, grid_285}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_286 = {{1'd0}, grid_286}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_287 = {{1'd0}, grid_287}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_288 = {{1'd0}, grid_288}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_289 = {{1'd0}, grid_289}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_290 = {{1'd0}, grid_290}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_291 = {{1'd0}, grid_291}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_292 = {{1'd0}, grid_292}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_293 = {{1'd0}, grid_293}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_294 = {{1'd0}, grid_294}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_295 = {{1'd0}, grid_295}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_296 = {{1'd0}, grid_296}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_297 = {{1'd0}, grid_297}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_298 = {{1'd0}, grid_298}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_grid_299 = {{1'd0}, grid_299}; // @[\\src\\main\\scala\\GameLogic.scala 113:28]
  assign movementDetector_io_xPos = 2'h0 == stateReg ? $signed(blockXReg) : $signed(_GEN_3130); // @[\\src\\main\\scala\\GameLogic.scala 186:20 114:28]
  assign movementDetector_io_yPos = 2'h0 == stateReg ? $signed(blockYReg) : $signed(_GEN_3133); // @[\\src\\main\\scala\\GameLogic.scala 186:20 115:28]
  assign movementDetector_io_xOffsets_0 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3143); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  assign movementDetector_io_xOffsets_1 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3144); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  assign movementDetector_io_xOffsets_2 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3145); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  assign movementDetector_io_xOffsets_3 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3146); // @[\\src\\main\\scala\\GameLogic.scala 186:20 116:32]
  assign movementDetector_io_yOffsets_0 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3147); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  assign movementDetector_io_yOffsets_1 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3148); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  assign movementDetector_io_yOffsets_2 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3149); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  assign movementDetector_io_yOffsets_3 = 2'h0 == stateReg ? $signed(4'sh0) : $signed(_GEN_3150); // @[\\src\\main\\scala\\GameLogic.scala 186:20 117:32]
  assign posToIndex_io_xPos = 2'h0 == stateReg ? $signed(11'sh0) : $signed(_GEN_2813); // @[\\src\\main\\scala\\GameLogic.scala 186:20 121:22]
  assign posToIndex_io_yPos = 2'h0 == stateReg ? $signed(10'sh0) : $signed(_GEN_2814); // @[\\src\\main\\scala\\GameLogic.scala 186:20 122:22]
  assign posToGridIndex_io_xPos = 2'h0 == stateReg ? $signed(11'sh0) : $signed(_GEN_2813); // @[\\src\\main\\scala\\GameLogic.scala 186:20 124:26]
  assign posToGridIndex_io_yPos = 2'h0 == stateReg ? $signed(10'sh0) : $signed(_GEN_2814); // @[\\src\\main\\scala\\GameLogic.scala 186:20 125:26]
  assign gameScreen_clock = clock;
  assign gameScreen_reset = reset;
  assign gameScreen_io_sw = io_sw_7; // @[\\src\\main\\scala\\GameLogic.scala 152:20]
  assign blockType_prng_clock = clock;
  assign blockType_prng_reset = reset;
  assign blockType_prng_io_increment = 1'h1; // @[src/main/scala/chisel3/util/random/PRNG.scala 94:23]
  assign rnd_prng_clock = clock;
  assign rnd_prng_reset = reset;
  assign rnd_prng_io_increment = 2'h0 == stateReg ? 1'h0 : _GEN_3127; // @[\\src\\main\\scala\\GameLogic.scala 186:20 193:17]
  assign blockLogic_io_rotation = rotation; // @[\\src\\main\\scala\\GameLogic.scala 170:26]
  assign blockLogic_io_xPos = blockXReg; // @[\\src\\main\\scala\\GameLogic.scala 168:22]
  assign blockLogic_io_yPos = blockYReg; // @[\\src\\main\\scala\\GameLogic.scala 169:22]
  assign blockLogic_io_sel = blockType; // @[\\src\\main\\scala\\GameLogic.scala 171:21]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 80:28]
      currentTask <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 80:28]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          currentTask <= _GEN_313;
        end
      end else if (2'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        currentTask <= _GEN_2770;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 81:29]
      writingCount <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 81:29]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          writingCount <= _GEN_310;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 84:29]
      currentBlock <= 4'h0; // @[\\src\\main\\scala\\GameLogic.scala 84:29]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (!(2'h1 == currentTask)) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          currentBlock <= _GEN_2133;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_0 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_0 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_0 <= _GEN_10;
      end else begin
        grid_0 <= _GEN_2136;
      end
    end else begin
      grid_0 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_1 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_1 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_1 <= _GEN_11;
      end else begin
        grid_1 <= _GEN_2137;
      end
    end else begin
      grid_1 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_2 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_2 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_2 <= _GEN_12;
      end else begin
        grid_2 <= _GEN_2138;
      end
    end else begin
      grid_2 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_3 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_3 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_3 <= _GEN_13;
      end else begin
        grid_3 <= _GEN_2139;
      end
    end else begin
      grid_3 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_4 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_4 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_4 <= _GEN_14;
      end else begin
        grid_4 <= _GEN_2140;
      end
    end else begin
      grid_4 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_5 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_5 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_5 <= _GEN_15;
      end else begin
        grid_5 <= _GEN_2141;
      end
    end else begin
      grid_5 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_6 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_6 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_6 <= _GEN_16;
      end else begin
        grid_6 <= _GEN_2142;
      end
    end else begin
      grid_6 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_7 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_7 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_7 <= _GEN_17;
      end else begin
        grid_7 <= _GEN_2143;
      end
    end else begin
      grid_7 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_8 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_8 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_8 <= _GEN_18;
      end else begin
        grid_8 <= _GEN_2144;
      end
    end else begin
      grid_8 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_9 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_9 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_9 <= _GEN_19;
      end else begin
        grid_9 <= _GEN_2145;
      end
    end else begin
      grid_9 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_10 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_10 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_10 <= _GEN_20;
      end else begin
        grid_10 <= _GEN_2146;
      end
    end else begin
      grid_10 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_11 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_11 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_11 <= _GEN_21;
      end else begin
        grid_11 <= _GEN_2147;
      end
    end else begin
      grid_11 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_12 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_12 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_12 <= _GEN_22;
      end else begin
        grid_12 <= _GEN_2148;
      end
    end else begin
      grid_12 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_13 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_13 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_13 <= _GEN_23;
      end else begin
        grid_13 <= _GEN_2149;
      end
    end else begin
      grid_13 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_14 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_14 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_14 <= _GEN_24;
      end else begin
        grid_14 <= _GEN_2150;
      end
    end else begin
      grid_14 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_15 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_15 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_15 <= _GEN_25;
      end else begin
        grid_15 <= _GEN_2151;
      end
    end else begin
      grid_15 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_16 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_16 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_16 <= _GEN_26;
      end else begin
        grid_16 <= _GEN_2152;
      end
    end else begin
      grid_16 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_17 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_17 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_17 <= _GEN_27;
      end else begin
        grid_17 <= _GEN_2153;
      end
    end else begin
      grid_17 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_18 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_18 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_18 <= _GEN_28;
      end else begin
        grid_18 <= _GEN_2154;
      end
    end else begin
      grid_18 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_19 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_19 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_19 <= _GEN_29;
      end else begin
        grid_19 <= _GEN_2155;
      end
    end else begin
      grid_19 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_20 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_20 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_20 <= _GEN_30;
      end else begin
        grid_20 <= _GEN_2156;
      end
    end else begin
      grid_20 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_21 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_21 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_21 <= _GEN_31;
      end else begin
        grid_21 <= _GEN_2157;
      end
    end else begin
      grid_21 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_22 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_22 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_22 <= _GEN_32;
      end else begin
        grid_22 <= _GEN_2158;
      end
    end else begin
      grid_22 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_23 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_23 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_23 <= _GEN_33;
      end else begin
        grid_23 <= _GEN_2159;
      end
    end else begin
      grid_23 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_24 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_24 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_24 <= _GEN_34;
      end else begin
        grid_24 <= _GEN_2160;
      end
    end else begin
      grid_24 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 95:13]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_25 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_25 <= _GEN_35;
        end else begin
          grid_25 <= _GEN_2161;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_26 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_26 <= _GEN_36;
        end else begin
          grid_26 <= _GEN_2162;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_27 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_27 <= _GEN_37;
        end else begin
          grid_27 <= _GEN_2163;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_28 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_28 <= _GEN_38;
        end else begin
          grid_28 <= _GEN_2164;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_29 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_29 <= _GEN_39;
        end else begin
          grid_29 <= _GEN_2165;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_30 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_30 <= _GEN_40;
        end else begin
          grid_30 <= _GEN_2166;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_31 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_31 <= _GEN_41;
        end else begin
          grid_31 <= _GEN_2167;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_32 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_32 <= _GEN_42;
        end else begin
          grid_32 <= _GEN_2168;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_33 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_33 <= _GEN_43;
        end else begin
          grid_33 <= _GEN_2169;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_34 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_34 <= _GEN_44;
        end else begin
          grid_34 <= _GEN_2170;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_35 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_35 <= _GEN_45;
        end else begin
          grid_35 <= _GEN_2171;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_36 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_36 <= _GEN_46;
        end else begin
          grid_36 <= _GEN_2172;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_37 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_37 <= _GEN_47;
        end else begin
          grid_37 <= _GEN_2173;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_38 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_38 <= _GEN_48;
        end else begin
          grid_38 <= _GEN_2174;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_39 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_39 <= _GEN_49;
        end else begin
          grid_39 <= _GEN_2175;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_40 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_40 <= _GEN_50;
        end else begin
          grid_40 <= _GEN_2176;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_41 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_41 <= _GEN_51;
        end else begin
          grid_41 <= _GEN_2177;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_42 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_42 <= _GEN_52;
        end else begin
          grid_42 <= _GEN_2178;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_43 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_43 <= _GEN_53;
        end else begin
          grid_43 <= _GEN_2179;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_44 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_44 <= _GEN_54;
        end else begin
          grid_44 <= _GEN_2180;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_45 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_45 <= _GEN_55;
        end else begin
          grid_45 <= _GEN_2181;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_46 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_46 <= _GEN_56;
        end else begin
          grid_46 <= _GEN_2182;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_47 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_47 <= _GEN_57;
        end else begin
          grid_47 <= _GEN_2183;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_48 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_48 <= _GEN_58;
        end else begin
          grid_48 <= _GEN_2184;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_49 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_49 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_49 <= _GEN_59;
      end else begin
        grid_49 <= _GEN_2185;
      end
    end else begin
      grid_49 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_50 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_50 <= _GEN_60;
        end else begin
          grid_50 <= _GEN_2186;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_51 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_51 <= _GEN_61;
        end else begin
          grid_51 <= _GEN_2187;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_52 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_52 <= _GEN_62;
        end else begin
          grid_52 <= _GEN_2188;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_53 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_53 <= _GEN_63;
        end else begin
          grid_53 <= _GEN_2189;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_54 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_54 <= _GEN_64;
        end else begin
          grid_54 <= _GEN_2190;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_55 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_55 <= _GEN_65;
        end else begin
          grid_55 <= _GEN_2191;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_56 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_56 <= _GEN_66;
        end else begin
          grid_56 <= _GEN_2192;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_57 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_57 <= _GEN_67;
        end else begin
          grid_57 <= _GEN_2193;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_58 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_58 <= _GEN_68;
        end else begin
          grid_58 <= _GEN_2194;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_59 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_59 <= _GEN_69;
        end else begin
          grid_59 <= _GEN_2195;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_60 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_60 <= _GEN_70;
        end else begin
          grid_60 <= _GEN_2196;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_61 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_61 <= _GEN_71;
        end else begin
          grid_61 <= _GEN_2197;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_62 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_62 <= _GEN_72;
        end else begin
          grid_62 <= _GEN_2198;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_63 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_63 <= _GEN_73;
        end else begin
          grid_63 <= _GEN_2199;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_64 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_64 <= _GEN_74;
        end else begin
          grid_64 <= _GEN_2200;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_65 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_65 <= _GEN_75;
        end else begin
          grid_65 <= _GEN_2201;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_66 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_66 <= _GEN_76;
        end else begin
          grid_66 <= _GEN_2202;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_67 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_67 <= _GEN_77;
        end else begin
          grid_67 <= _GEN_2203;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_68 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_68 <= _GEN_78;
        end else begin
          grid_68 <= _GEN_2204;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_69 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_69 <= _GEN_79;
        end else begin
          grid_69 <= _GEN_2205;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_70 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_70 <= _GEN_80;
        end else begin
          grid_70 <= _GEN_2206;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_71 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_71 <= _GEN_81;
        end else begin
          grid_71 <= _GEN_2207;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_72 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_72 <= _GEN_82;
        end else begin
          grid_72 <= _GEN_2208;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_73 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_73 <= _GEN_83;
        end else begin
          grid_73 <= _GEN_2209;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_74 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_74 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_74 <= _GEN_84;
      end else begin
        grid_74 <= _GEN_2210;
      end
    end else begin
      grid_74 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_75 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_75 <= _GEN_85;
        end else begin
          grid_75 <= _GEN_2211;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_76 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_76 <= _GEN_86;
        end else begin
          grid_76 <= _GEN_2212;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_77 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_77 <= _GEN_87;
        end else begin
          grid_77 <= _GEN_2213;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_78 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_78 <= _GEN_88;
        end else begin
          grid_78 <= _GEN_2214;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_79 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_79 <= _GEN_89;
        end else begin
          grid_79 <= _GEN_2215;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_80 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_80 <= _GEN_90;
        end else begin
          grid_80 <= _GEN_2216;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_81 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_81 <= _GEN_91;
        end else begin
          grid_81 <= _GEN_2217;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_82 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_82 <= _GEN_92;
        end else begin
          grid_82 <= _GEN_2218;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_83 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_83 <= _GEN_93;
        end else begin
          grid_83 <= _GEN_2219;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_84 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_84 <= _GEN_94;
        end else begin
          grid_84 <= _GEN_2220;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_85 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_85 <= _GEN_95;
        end else begin
          grid_85 <= _GEN_2221;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_86 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_86 <= _GEN_96;
        end else begin
          grid_86 <= _GEN_2222;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_87 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_87 <= _GEN_97;
        end else begin
          grid_87 <= _GEN_2223;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_88 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_88 <= _GEN_98;
        end else begin
          grid_88 <= _GEN_2224;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_89 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_89 <= _GEN_99;
        end else begin
          grid_89 <= _GEN_2225;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_90 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_90 <= _GEN_100;
        end else begin
          grid_90 <= _GEN_2226;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_91 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_91 <= _GEN_101;
        end else begin
          grid_91 <= _GEN_2227;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_92 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_92 <= _GEN_102;
        end else begin
          grid_92 <= _GEN_2228;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_93 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_93 <= _GEN_103;
        end else begin
          grid_93 <= _GEN_2229;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_94 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_94 <= _GEN_104;
        end else begin
          grid_94 <= _GEN_2230;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_95 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_95 <= _GEN_105;
        end else begin
          grid_95 <= _GEN_2231;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_96 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_96 <= _GEN_106;
        end else begin
          grid_96 <= _GEN_2232;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_97 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_97 <= _GEN_107;
        end else begin
          grid_97 <= _GEN_2233;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_98 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_98 <= _GEN_108;
        end else begin
          grid_98 <= _GEN_2234;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_99 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_99 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_99 <= _GEN_109;
      end else begin
        grid_99 <= _GEN_2235;
      end
    end else begin
      grid_99 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_100 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_100 <= _GEN_110;
        end else begin
          grid_100 <= _GEN_2236;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_101 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_101 <= _GEN_111;
        end else begin
          grid_101 <= _GEN_2237;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_102 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_102 <= _GEN_112;
        end else begin
          grid_102 <= _GEN_2238;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_103 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_103 <= _GEN_113;
        end else begin
          grid_103 <= _GEN_2239;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_104 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_104 <= _GEN_114;
        end else begin
          grid_104 <= _GEN_2240;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_105 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_105 <= _GEN_115;
        end else begin
          grid_105 <= _GEN_2241;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_106 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_106 <= _GEN_116;
        end else begin
          grid_106 <= _GEN_2242;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_107 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_107 <= _GEN_117;
        end else begin
          grid_107 <= _GEN_2243;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_108 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_108 <= _GEN_118;
        end else begin
          grid_108 <= _GEN_2244;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_109 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_109 <= _GEN_119;
        end else begin
          grid_109 <= _GEN_2245;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_110 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_110 <= _GEN_120;
        end else begin
          grid_110 <= _GEN_2246;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_111 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_111 <= _GEN_121;
        end else begin
          grid_111 <= _GEN_2247;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_112 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_112 <= _GEN_122;
        end else begin
          grid_112 <= _GEN_2248;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_113 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_113 <= _GEN_123;
        end else begin
          grid_113 <= _GEN_2249;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_114 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_114 <= _GEN_124;
        end else begin
          grid_114 <= _GEN_2250;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_115 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_115 <= _GEN_125;
        end else begin
          grid_115 <= _GEN_2251;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_116 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_116 <= _GEN_126;
        end else begin
          grid_116 <= _GEN_2252;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_117 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_117 <= _GEN_127;
        end else begin
          grid_117 <= _GEN_2253;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_118 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_118 <= _GEN_128;
        end else begin
          grid_118 <= _GEN_2254;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_119 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_119 <= _GEN_129;
        end else begin
          grid_119 <= _GEN_2255;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_120 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_120 <= _GEN_130;
        end else begin
          grid_120 <= _GEN_2256;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_121 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_121 <= _GEN_131;
        end else begin
          grid_121 <= _GEN_2257;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_122 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_122 <= _GEN_132;
        end else begin
          grid_122 <= _GEN_2258;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_123 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_123 <= _GEN_133;
        end else begin
          grid_123 <= _GEN_2259;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_124 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_124 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_124 <= _GEN_134;
      end else begin
        grid_124 <= _GEN_2260;
      end
    end else begin
      grid_124 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_125 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_125 <= _GEN_135;
        end else begin
          grid_125 <= _GEN_2261;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_126 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_126 <= _GEN_136;
        end else begin
          grid_126 <= _GEN_2262;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_127 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_127 <= _GEN_137;
        end else begin
          grid_127 <= _GEN_2263;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_128 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_128 <= _GEN_138;
        end else begin
          grid_128 <= _GEN_2264;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_129 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_129 <= _GEN_139;
        end else begin
          grid_129 <= _GEN_2265;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_130 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_130 <= _GEN_140;
        end else begin
          grid_130 <= _GEN_2266;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_131 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_131 <= _GEN_141;
        end else begin
          grid_131 <= _GEN_2267;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_132 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_132 <= _GEN_142;
        end else begin
          grid_132 <= _GEN_2268;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_133 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_133 <= _GEN_143;
        end else begin
          grid_133 <= _GEN_2269;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_134 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_134 <= _GEN_144;
        end else begin
          grid_134 <= _GEN_2270;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_135 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_135 <= _GEN_145;
        end else begin
          grid_135 <= _GEN_2271;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_136 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_136 <= _GEN_146;
        end else begin
          grid_136 <= _GEN_2272;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_137 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_137 <= _GEN_147;
        end else begin
          grid_137 <= _GEN_2273;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_138 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_138 <= _GEN_148;
        end else begin
          grid_138 <= _GEN_2274;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_139 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_139 <= _GEN_149;
        end else begin
          grid_139 <= _GEN_2275;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_140 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_140 <= _GEN_150;
        end else begin
          grid_140 <= _GEN_2276;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_141 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_141 <= _GEN_151;
        end else begin
          grid_141 <= _GEN_2277;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_142 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_142 <= _GEN_152;
        end else begin
          grid_142 <= _GEN_2278;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_143 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_143 <= _GEN_153;
        end else begin
          grid_143 <= _GEN_2279;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_144 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_144 <= _GEN_154;
        end else begin
          grid_144 <= _GEN_2280;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_145 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_145 <= _GEN_155;
        end else begin
          grid_145 <= _GEN_2281;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_146 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_146 <= _GEN_156;
        end else begin
          grid_146 <= _GEN_2282;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_147 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_147 <= _GEN_157;
        end else begin
          grid_147 <= _GEN_2283;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_148 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_148 <= _GEN_158;
        end else begin
          grid_148 <= _GEN_2284;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_149 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_149 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_149 <= _GEN_159;
      end else begin
        grid_149 <= _GEN_2285;
      end
    end else begin
      grid_149 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_150 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_150 <= _GEN_160;
        end else begin
          grid_150 <= _GEN_2286;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_151 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_151 <= _GEN_161;
        end else begin
          grid_151 <= _GEN_2287;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_152 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_152 <= _GEN_162;
        end else begin
          grid_152 <= _GEN_2288;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_153 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_153 <= _GEN_163;
        end else begin
          grid_153 <= _GEN_2289;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_154 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_154 <= _GEN_164;
        end else begin
          grid_154 <= _GEN_2290;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_155 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_155 <= _GEN_165;
        end else begin
          grid_155 <= _GEN_2291;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_156 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_156 <= _GEN_166;
        end else begin
          grid_156 <= _GEN_2292;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_157 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_157 <= _GEN_167;
        end else begin
          grid_157 <= _GEN_2293;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_158 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_158 <= _GEN_168;
        end else begin
          grid_158 <= _GEN_2294;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_159 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_159 <= _GEN_169;
        end else begin
          grid_159 <= _GEN_2295;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_160 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_160 <= _GEN_170;
        end else begin
          grid_160 <= _GEN_2296;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_161 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_161 <= _GEN_171;
        end else begin
          grid_161 <= _GEN_2297;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_162 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_162 <= _GEN_172;
        end else begin
          grid_162 <= _GEN_2298;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_163 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_163 <= _GEN_173;
        end else begin
          grid_163 <= _GEN_2299;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_164 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_164 <= _GEN_174;
        end else begin
          grid_164 <= _GEN_2300;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_165 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_165 <= _GEN_175;
        end else begin
          grid_165 <= _GEN_2301;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_166 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_166 <= _GEN_176;
        end else begin
          grid_166 <= _GEN_2302;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_167 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_167 <= _GEN_177;
        end else begin
          grid_167 <= _GEN_2303;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_168 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_168 <= _GEN_178;
        end else begin
          grid_168 <= _GEN_2304;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_169 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_169 <= _GEN_179;
        end else begin
          grid_169 <= _GEN_2305;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_170 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_170 <= _GEN_180;
        end else begin
          grid_170 <= _GEN_2306;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_171 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_171 <= _GEN_181;
        end else begin
          grid_171 <= _GEN_2307;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_172 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_172 <= _GEN_182;
        end else begin
          grid_172 <= _GEN_2308;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_173 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_173 <= _GEN_183;
        end else begin
          grid_173 <= _GEN_2309;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_174 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_174 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_174 <= _GEN_184;
      end else begin
        grid_174 <= _GEN_2310;
      end
    end else begin
      grid_174 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_175 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_175 <= _GEN_185;
        end else begin
          grid_175 <= _GEN_2311;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_176 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_176 <= _GEN_186;
        end else begin
          grid_176 <= _GEN_2312;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_177 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_177 <= _GEN_187;
        end else begin
          grid_177 <= _GEN_2313;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_178 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_178 <= _GEN_188;
        end else begin
          grid_178 <= _GEN_2314;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_179 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_179 <= _GEN_189;
        end else begin
          grid_179 <= _GEN_2315;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_180 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_180 <= _GEN_190;
        end else begin
          grid_180 <= _GEN_2316;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_181 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_181 <= _GEN_191;
        end else begin
          grid_181 <= _GEN_2317;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_182 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_182 <= _GEN_192;
        end else begin
          grid_182 <= _GEN_2318;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_183 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_183 <= _GEN_193;
        end else begin
          grid_183 <= _GEN_2319;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_184 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_184 <= _GEN_194;
        end else begin
          grid_184 <= _GEN_2320;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_185 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_185 <= _GEN_195;
        end else begin
          grid_185 <= _GEN_2321;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_186 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_186 <= _GEN_196;
        end else begin
          grid_186 <= _GEN_2322;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_187 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_187 <= _GEN_197;
        end else begin
          grid_187 <= _GEN_2323;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_188 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_188 <= _GEN_198;
        end else begin
          grid_188 <= _GEN_2324;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_189 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_189 <= _GEN_199;
        end else begin
          grid_189 <= _GEN_2325;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_190 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_190 <= _GEN_200;
        end else begin
          grid_190 <= _GEN_2326;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_191 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_191 <= _GEN_201;
        end else begin
          grid_191 <= _GEN_2327;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_192 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_192 <= _GEN_202;
        end else begin
          grid_192 <= _GEN_2328;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_193 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_193 <= _GEN_203;
        end else begin
          grid_193 <= _GEN_2329;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_194 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_194 <= _GEN_204;
        end else begin
          grid_194 <= _GEN_2330;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_195 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_195 <= _GEN_205;
        end else begin
          grid_195 <= _GEN_2331;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_196 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_196 <= _GEN_206;
        end else begin
          grid_196 <= _GEN_2332;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_197 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_197 <= _GEN_207;
        end else begin
          grid_197 <= _GEN_2333;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_198 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_198 <= _GEN_208;
        end else begin
          grid_198 <= _GEN_2334;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_199 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_199 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_199 <= _GEN_209;
      end else begin
        grid_199 <= _GEN_2335;
      end
    end else begin
      grid_199 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_200 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_200 <= _GEN_210;
        end else begin
          grid_200 <= _GEN_2336;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_201 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_201 <= _GEN_211;
        end else begin
          grid_201 <= _GEN_2337;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_202 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_202 <= _GEN_212;
        end else begin
          grid_202 <= _GEN_2338;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_203 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_203 <= _GEN_213;
        end else begin
          grid_203 <= _GEN_2339;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_204 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_204 <= _GEN_214;
        end else begin
          grid_204 <= _GEN_2340;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_205 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_205 <= _GEN_215;
        end else begin
          grid_205 <= _GEN_2341;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_206 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_206 <= _GEN_216;
        end else begin
          grid_206 <= _GEN_2342;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_207 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_207 <= _GEN_217;
        end else begin
          grid_207 <= _GEN_2343;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_208 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_208 <= _GEN_218;
        end else begin
          grid_208 <= _GEN_2344;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_209 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_209 <= _GEN_219;
        end else begin
          grid_209 <= _GEN_2345;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_210 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_210 <= _GEN_220;
        end else begin
          grid_210 <= _GEN_2346;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_211 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_211 <= _GEN_221;
        end else begin
          grid_211 <= _GEN_2347;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_212 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_212 <= _GEN_222;
        end else begin
          grid_212 <= _GEN_2348;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_213 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_213 <= _GEN_223;
        end else begin
          grid_213 <= _GEN_2349;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_214 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_214 <= _GEN_224;
        end else begin
          grid_214 <= _GEN_2350;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_215 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_215 <= _GEN_225;
        end else begin
          grid_215 <= _GEN_2351;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_216 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_216 <= _GEN_226;
        end else begin
          grid_216 <= _GEN_2352;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_217 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_217 <= _GEN_227;
        end else begin
          grid_217 <= _GEN_2353;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_218 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_218 <= _GEN_228;
        end else begin
          grid_218 <= _GEN_2354;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_219 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_219 <= _GEN_229;
        end else begin
          grid_219 <= _GEN_2355;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_220 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_220 <= _GEN_230;
        end else begin
          grid_220 <= _GEN_2356;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_221 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_221 <= _GEN_231;
        end else begin
          grid_221 <= _GEN_2357;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_222 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_222 <= _GEN_232;
        end else begin
          grid_222 <= _GEN_2358;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_223 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_223 <= _GEN_233;
        end else begin
          grid_223 <= _GEN_2359;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_224 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_224 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_224 <= _GEN_234;
      end else begin
        grid_224 <= _GEN_2360;
      end
    end else begin
      grid_224 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_225 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_225 <= _GEN_235;
        end else begin
          grid_225 <= _GEN_2361;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_226 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_226 <= _GEN_236;
        end else begin
          grid_226 <= _GEN_2362;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_227 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_227 <= _GEN_237;
        end else begin
          grid_227 <= _GEN_2363;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_228 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_228 <= _GEN_238;
        end else begin
          grid_228 <= _GEN_2364;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_229 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_229 <= _GEN_239;
        end else begin
          grid_229 <= _GEN_2365;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_230 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_230 <= _GEN_240;
        end else begin
          grid_230 <= _GEN_2366;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_231 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_231 <= _GEN_241;
        end else begin
          grid_231 <= _GEN_2367;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_232 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_232 <= _GEN_242;
        end else begin
          grid_232 <= _GEN_2368;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_233 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_233 <= _GEN_243;
        end else begin
          grid_233 <= _GEN_2369;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_234 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_234 <= _GEN_244;
        end else begin
          grid_234 <= _GEN_2370;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_235 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_235 <= _GEN_245;
        end else begin
          grid_235 <= _GEN_2371;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_236 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_236 <= _GEN_246;
        end else begin
          grid_236 <= _GEN_2372;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_237 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_237 <= _GEN_247;
        end else begin
          grid_237 <= _GEN_2373;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_238 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_238 <= _GEN_248;
        end else begin
          grid_238 <= _GEN_2374;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_239 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_239 <= _GEN_249;
        end else begin
          grid_239 <= _GEN_2375;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_240 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_240 <= _GEN_250;
        end else begin
          grid_240 <= _GEN_2376;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_241 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_241 <= _GEN_251;
        end else begin
          grid_241 <= _GEN_2377;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_242 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_242 <= _GEN_252;
        end else begin
          grid_242 <= _GEN_2378;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_243 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_243 <= _GEN_253;
        end else begin
          grid_243 <= _GEN_2379;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_244 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_244 <= _GEN_254;
        end else begin
          grid_244 <= _GEN_2380;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_245 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_245 <= _GEN_255;
        end else begin
          grid_245 <= _GEN_2381;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_246 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_246 <= _GEN_256;
        end else begin
          grid_246 <= _GEN_2382;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_247 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_247 <= _GEN_257;
        end else begin
          grid_247 <= _GEN_2383;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_248 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_248 <= _GEN_258;
        end else begin
          grid_248 <= _GEN_2384;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_249 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_249 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_249 <= _GEN_259;
      end else begin
        grid_249 <= _GEN_2385;
      end
    end else begin
      grid_249 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_250 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_250 <= _GEN_260;
        end else begin
          grid_250 <= _GEN_2386;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_251 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_251 <= _GEN_261;
        end else begin
          grid_251 <= _GEN_2387;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_252 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_252 <= _GEN_262;
        end else begin
          grid_252 <= _GEN_2388;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_253 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_253 <= _GEN_263;
        end else begin
          grid_253 <= _GEN_2389;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_254 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_254 <= _GEN_264;
        end else begin
          grid_254 <= _GEN_2390;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_255 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_255 <= _GEN_265;
        end else begin
          grid_255 <= _GEN_2391;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_256 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_256 <= _GEN_266;
        end else begin
          grid_256 <= _GEN_2392;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_257 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_257 <= _GEN_267;
        end else begin
          grid_257 <= _GEN_2393;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_258 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_258 <= _GEN_268;
        end else begin
          grid_258 <= _GEN_2394;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_259 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_259 <= _GEN_269;
        end else begin
          grid_259 <= _GEN_2395;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_260 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_260 <= _GEN_270;
        end else begin
          grid_260 <= _GEN_2396;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_261 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_261 <= _GEN_271;
        end else begin
          grid_261 <= _GEN_2397;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_262 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_262 <= _GEN_272;
        end else begin
          grid_262 <= _GEN_2398;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_263 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_263 <= _GEN_273;
        end else begin
          grid_263 <= _GEN_2399;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_264 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_264 <= _GEN_274;
        end else begin
          grid_264 <= _GEN_2400;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_265 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_265 <= _GEN_275;
        end else begin
          grid_265 <= _GEN_2401;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_266 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_266 <= _GEN_276;
        end else begin
          grid_266 <= _GEN_2402;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_267 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_267 <= _GEN_277;
        end else begin
          grid_267 <= _GEN_2403;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_268 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_268 <= _GEN_278;
        end else begin
          grid_268 <= _GEN_2404;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_269 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_269 <= _GEN_279;
        end else begin
          grid_269 <= _GEN_2405;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_270 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_270 <= _GEN_280;
        end else begin
          grid_270 <= _GEN_2406;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_271 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_271 <= _GEN_281;
        end else begin
          grid_271 <= _GEN_2407;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_272 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_272 <= _GEN_282;
        end else begin
          grid_272 <= _GEN_2408;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_273 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          grid_273 <= _GEN_283;
        end else begin
          grid_273 <= _GEN_2409;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_274 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_274 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_274 <= _GEN_284;
      end else begin
        grid_274 <= _GEN_2410;
      end
    end else begin
      grid_274 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 91:23]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_275 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_275 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_275 <= _GEN_285;
      end else begin
        grid_275 <= _GEN_2411;
      end
    end else begin
      grid_275 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_276 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_276 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_276 <= _GEN_286;
      end else begin
        grid_276 <= _GEN_2412;
      end
    end else begin
      grid_276 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_277 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_277 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_277 <= _GEN_287;
      end else begin
        grid_277 <= _GEN_2413;
      end
    end else begin
      grid_277 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_278 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_278 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_278 <= _GEN_288;
      end else begin
        grid_278 <= _GEN_2414;
      end
    end else begin
      grid_278 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_279 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_279 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_279 <= _GEN_289;
      end else begin
        grid_279 <= _GEN_2415;
      end
    end else begin
      grid_279 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_280 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_280 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_280 <= _GEN_290;
      end else begin
        grid_280 <= _GEN_2416;
      end
    end else begin
      grid_280 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_281 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_281 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_281 <= _GEN_291;
      end else begin
        grid_281 <= _GEN_2417;
      end
    end else begin
      grid_281 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_282 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_282 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_282 <= _GEN_292;
      end else begin
        grid_282 <= _GEN_2418;
      end
    end else begin
      grid_282 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_283 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_283 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_283 <= _GEN_293;
      end else begin
        grid_283 <= _GEN_2419;
      end
    end else begin
      grid_283 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_284 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_284 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_284 <= _GEN_294;
      end else begin
        grid_284 <= _GEN_2420;
      end
    end else begin
      grid_284 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_285 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_285 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_285 <= _GEN_295;
      end else begin
        grid_285 <= _GEN_2421;
      end
    end else begin
      grid_285 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_286 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_286 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_286 <= _GEN_296;
      end else begin
        grid_286 <= _GEN_2422;
      end
    end else begin
      grid_286 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_287 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_287 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_287 <= _GEN_297;
      end else begin
        grid_287 <= _GEN_2423;
      end
    end else begin
      grid_287 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_288 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_288 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_288 <= _GEN_298;
      end else begin
        grid_288 <= _GEN_2424;
      end
    end else begin
      grid_288 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_289 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_289 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_289 <= _GEN_299;
      end else begin
        grid_289 <= _GEN_2425;
      end
    end else begin
      grid_289 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_290 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_290 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_290 <= _GEN_300;
      end else begin
        grid_290 <= _GEN_2426;
      end
    end else begin
      grid_290 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_291 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_291 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_291 <= _GEN_301;
      end else begin
        grid_291 <= _GEN_2427;
      end
    end else begin
      grid_291 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_292 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_292 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_292 <= _GEN_302;
      end else begin
        grid_292 <= _GEN_2428;
      end
    end else begin
      grid_292 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_293 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_293 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_293 <= _GEN_303;
      end else begin
        grid_293 <= _GEN_2429;
      end
    end else begin
      grid_293 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_294 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_294 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_294 <= _GEN_304;
      end else begin
        grid_294 <= _GEN_2430;
      end
    end else begin
      grid_294 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_295 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_295 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_295 <= _GEN_305;
      end else begin
        grid_295 <= _GEN_2431;
      end
    end else begin
      grid_295 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_296 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_296 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_296 <= _GEN_306;
      end else begin
        grid_296 <= _GEN_2432;
      end
    end else begin
      grid_296 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_297 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_297 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_297 <= _GEN_307;
      end else begin
        grid_297 <= _GEN_2433;
      end
    end else begin
      grid_297 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_298 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_298 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_298 <= _GEN_308;
      end else begin
        grid_298 <= _GEN_2434;
      end
    end else begin
      grid_298 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 88:21]
      grid_299 <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 88:21]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      grid_299 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        grid_299 <= _GEN_309;
      end else begin
        grid_299 <= _GEN_2435;
      end
    end else begin
      grid_299 <= 2'h1; // @[\\src\\main\\scala\\GameLogic.scala 96:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 102:26]
      blockXReg <= -11'sh4; // @[\\src\\main\\scala\\GameLogic.scala 102:26]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          blockXReg <= _GEN_311;
        end
      end else if (2'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        blockXReg <= _GEN_2765;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 103:26]
      blockYReg <= 10'sh8; // @[\\src\\main\\scala\\GameLogic.scala 103:26]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          blockYReg <= _GEN_312;
        end
      end else if (2'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        blockYReg <= _GEN_2766;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 137:25]
      stateReg <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 137:25]
    end else if (2'h0 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (io_newFrame & ~gameScreen_io_staticScreen) begin // @[\\src\\main\\scala\\GameLogic.scala 188:56]
        stateReg <= 2'h2; // @[\\src\\main\\scala\\GameLogic.scala 189:18]
      end else if (gameScreen_io_staticScreen) begin // @[\\src\\main\\scala\\GameLogic.scala 190:47]
        stateReg <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 191:18]
      end
    end else if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
        stateReg <= _GEN_314;
      end else begin
        stateReg <= _GEN_2132;
      end
    end else if (2'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      stateReg <= nextState; // @[\\src\\main\\scala\\GameLogic.scala 315:16]
    end else begin
      stateReg <= _GEN_2780;
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 142:24]
      moveCnt <= 7'h0; // @[\\src\\main\\scala\\GameLogic.scala 142:24]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (!(2'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
          moveCnt <= _GEN_2753;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 147:25]
      rotation <= 2'h0; // @[\\src\\main\\scala\\GameLogic.scala 147:25]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          rotation <= _GEN_316;
        end
      end else if (2'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        rotation <= _GEN_2767;
      end
    end
    upRelease <= reset | _GEN_3474; // @[\\src\\main\\scala\\GameLogic.scala 149:{26,26}]
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 157:26]
      blockType <= _blockType_T; // @[\\src\\main\\scala\\GameLogic.scala 157:26]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (!(2'h1 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
          blockType <= _GEN_2751;
        end
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 165:25]
      newPiece <= 1'h0; // @[\\src\\main\\scala\\GameLogic.scala 165:25]
    end else if (!(2'h0 == stateReg)) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
      if (2'h1 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        if (2'h1 == currentTask) begin // @[\\src\\main\\scala\\GameLogic.scala 196:27]
          newPiece <= _GEN_315;
        end
      end else if (2'h2 == stateReg) begin // @[\\src\\main\\scala\\GameLogic.scala 186:20]
        newPiece <= _GEN_2752;
      end
    end
    if (reset) begin // @[\\src\\main\\scala\\GameLogic.scala 178:31]
      speedThreshold <= 7'h78; // @[\\src\\main\\scala\\GameLogic.scala 178:31]
    end else if (io_btnD) begin // @[\\src\\main\\scala\\GameLogic.scala 179:24]
      speedThreshold <= 7'h1e;
    end else begin
      speedThreshold <= 7'h78;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  currentTask = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  writingCount = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  currentBlock = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  grid_0 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  grid_1 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  grid_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  grid_3 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  grid_4 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  grid_5 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  grid_6 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  grid_7 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  grid_8 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  grid_9 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  grid_10 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  grid_11 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  grid_12 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  grid_13 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  grid_14 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  grid_15 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  grid_16 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  grid_17 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  grid_18 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  grid_19 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  grid_20 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  grid_21 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  grid_22 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  grid_23 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  grid_24 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  grid_25 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  grid_26 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  grid_27 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  grid_28 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  grid_29 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  grid_30 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  grid_31 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  grid_32 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  grid_33 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  grid_34 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  grid_35 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  grid_36 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  grid_37 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  grid_38 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  grid_39 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  grid_40 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  grid_41 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  grid_42 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  grid_43 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  grid_44 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  grid_45 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  grid_46 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  grid_47 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  grid_48 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  grid_49 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  grid_50 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  grid_51 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  grid_52 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  grid_53 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  grid_54 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  grid_55 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  grid_56 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  grid_57 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  grid_58 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  grid_59 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  grid_60 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  grid_61 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  grid_62 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  grid_63 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  grid_64 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  grid_65 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  grid_66 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  grid_67 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  grid_68 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  grid_69 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  grid_70 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  grid_71 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  grid_72 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  grid_73 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  grid_74 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  grid_75 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  grid_76 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  grid_77 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  grid_78 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  grid_79 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  grid_80 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  grid_81 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  grid_82 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  grid_83 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  grid_84 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  grid_85 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  grid_86 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  grid_87 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  grid_88 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  grid_89 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  grid_90 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  grid_91 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  grid_92 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  grid_93 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  grid_94 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  grid_95 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  grid_96 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  grid_97 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  grid_98 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  grid_99 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  grid_100 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  grid_101 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  grid_102 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  grid_103 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  grid_104 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  grid_105 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  grid_106 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  grid_107 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  grid_108 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  grid_109 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  grid_110 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  grid_111 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  grid_112 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  grid_113 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  grid_114 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  grid_115 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  grid_116 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  grid_117 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  grid_118 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  grid_119 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  grid_120 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  grid_121 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  grid_122 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  grid_123 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  grid_124 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  grid_125 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  grid_126 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  grid_127 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  grid_128 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  grid_129 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  grid_130 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  grid_131 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  grid_132 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  grid_133 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  grid_134 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  grid_135 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  grid_136 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  grid_137 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  grid_138 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  grid_139 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  grid_140 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  grid_141 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  grid_142 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  grid_143 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  grid_144 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  grid_145 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  grid_146 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  grid_147 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  grid_148 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  grid_149 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  grid_150 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  grid_151 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  grid_152 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  grid_153 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  grid_154 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  grid_155 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  grid_156 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  grid_157 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  grid_158 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  grid_159 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  grid_160 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  grid_161 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  grid_162 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  grid_163 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  grid_164 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  grid_165 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  grid_166 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  grid_167 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  grid_168 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  grid_169 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  grid_170 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  grid_171 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  grid_172 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  grid_173 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  grid_174 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  grid_175 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  grid_176 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  grid_177 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  grid_178 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  grid_179 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  grid_180 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  grid_181 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  grid_182 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  grid_183 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  grid_184 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  grid_185 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  grid_186 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  grid_187 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  grid_188 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  grid_189 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  grid_190 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  grid_191 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  grid_192 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  grid_193 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  grid_194 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  grid_195 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  grid_196 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  grid_197 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  grid_198 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  grid_199 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  grid_200 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  grid_201 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  grid_202 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  grid_203 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  grid_204 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  grid_205 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  grid_206 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  grid_207 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  grid_208 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  grid_209 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  grid_210 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  grid_211 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  grid_212 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  grid_213 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  grid_214 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  grid_215 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  grid_216 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  grid_217 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  grid_218 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  grid_219 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  grid_220 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  grid_221 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  grid_222 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  grid_223 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  grid_224 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  grid_225 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  grid_226 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  grid_227 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  grid_228 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  grid_229 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  grid_230 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  grid_231 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  grid_232 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  grid_233 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  grid_234 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  grid_235 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  grid_236 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  grid_237 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  grid_238 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  grid_239 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  grid_240 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  grid_241 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  grid_242 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  grid_243 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  grid_244 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  grid_245 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  grid_246 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  grid_247 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  grid_248 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  grid_249 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  grid_250 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  grid_251 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  grid_252 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  grid_253 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  grid_254 = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  grid_255 = _RAND_258[1:0];
  _RAND_259 = {1{`RANDOM}};
  grid_256 = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  grid_257 = _RAND_260[1:0];
  _RAND_261 = {1{`RANDOM}};
  grid_258 = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  grid_259 = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  grid_260 = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  grid_261 = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  grid_262 = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  grid_263 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  grid_264 = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  grid_265 = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  grid_266 = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  grid_267 = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  grid_268 = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  grid_269 = _RAND_272[1:0];
  _RAND_273 = {1{`RANDOM}};
  grid_270 = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  grid_271 = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  grid_272 = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  grid_273 = _RAND_276[1:0];
  _RAND_277 = {1{`RANDOM}};
  grid_274 = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  grid_275 = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  grid_276 = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  grid_277 = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  grid_278 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  grid_279 = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  grid_280 = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  grid_281 = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  grid_282 = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  grid_283 = _RAND_286[1:0];
  _RAND_287 = {1{`RANDOM}};
  grid_284 = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  grid_285 = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  grid_286 = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  grid_287 = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  grid_288 = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  grid_289 = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  grid_290 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  grid_291 = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  grid_292 = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  grid_293 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  grid_294 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  grid_295 = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  grid_296 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  grid_297 = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  grid_298 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  grid_299 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  blockXReg = _RAND_303[10:0];
  _RAND_304 = {1{`RANDOM}};
  blockYReg = _RAND_304[9:0];
  _RAND_305 = {1{`RANDOM}};
  stateReg = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  moveCnt = _RAND_306[6:0];
  _RAND_307 = {1{`RANDOM}};
  rotation = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  upRelease = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  blockType = _RAND_309[2:0];
  _RAND_310 = {1{`RANDOM}};
  newPiece = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  speedThreshold = _RAND_311[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GameTop(
  input        clock,
  input        reset,
  input        io_btnU, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnL, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnR, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_btnD, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaRed, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaBlue, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output [3:0] io_vgaGreen, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_Hsync, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_Vsync, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  input        io_sw_7, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_led_0, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_led_1, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_led_2, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_led_3, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_missingFrameError, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_backBufferWriteError, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_viewBoxOutOfRangeError, // @[\\src\\main\\scala\\GameTop.scala 14:14]
  output       io_soundOut // @[\\src\\main\\scala\\GameTop.scala 14:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  graphicEngineVGA_clock; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_reset; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_0; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_1; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_2; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_4; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_5; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_6; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_15; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_0; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_1; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_2; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_4; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_5; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_6; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_15; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_0; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_1; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_2; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [8:0] graphicEngineVGA_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [4:0] graphicEngineVGA_io_backBufferWriteData; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_backBufferWriteAddress; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_backBufferWriteEnable; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_missingFrameError; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_backBufferWriteError; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaRed; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaBlue; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaGreen; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Hsync; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Vsync; // @[\\src\\main\\scala\\GameTop.scala 46:32]
  wire  soundEngine_clock; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  soundEngine_reset; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  soundEngine_io_soundOut; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  soundEngine_io_startTune_0; // @[\\src\\main\\scala\\GameTop.scala 49:27]
  wire  gameLogic_clock; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_reset; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnU; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnL; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnR; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_btnD; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_sw_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_led_0; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_led_1; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_led_2; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_led_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_0; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_1; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_2; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_4; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_5; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_6; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_15; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_0; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_1; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_2; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_4; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_5; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_6; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_15; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_0; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_1; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_2; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [9:0] gameLogic_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [8:0] gameLogic_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [4:0] gameLogic_io_backBufferWriteData; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire [10:0] gameLogic_io_backBufferWriteAddress; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_backBufferWriteEnable; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  wire  gameLogic_io_startTune_0; // @[\\src\\main\\scala\\GameTop.scala 53:25]
  reg [20:0] debounceCounter; // @[\\src\\main\\scala\\GameTop.scala 59:32]
  wire  debounceSampleEn = debounceCounter == 21'h1e847f; // @[\\src\\main\\scala\\GameTop.scala 61:24]
  wire [20:0] _debounceCounter_T_1 = debounceCounter + 21'h1; // @[\\src\\main\\scala\\GameTop.scala 65:40]
  reg [21:0] resetReleaseCounter; // @[\\src\\main\\scala\\GameTop.scala 72:36]
  wire [21:0] _resetReleaseCounter_T_1 = resetReleaseCounter + 22'h1; // @[\\src\\main\\scala\\GameTop.scala 78:48]
  reg  btnUState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnUState; // @[\\src\\main\\scala\\GameTop.scala 85:28]
  reg  btnLState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnLState; // @[\\src\\main\\scala\\GameTop.scala 86:28]
  reg  btnRState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnRState; // @[\\src\\main\\scala\\GameTop.scala 87:28]
  reg  btnDState_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  btnDState; // @[\\src\\main\\scala\\GameTop.scala 88:28]
  reg  gameLogic_io_sw_7_pipeReg_0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  gameLogic_io_sw_7_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  gameLogic_io_sw_7_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
  reg  gameLogic_io_sw_7_r; // @[\\src\\main\\scala\\GameTop.scala 104:36]
  GraphicEngineVGA graphicEngineVGA ( // @[\\src\\main\\scala\\GameTop.scala 46:32]
    .clock(graphicEngineVGA_clock),
    .reset(graphicEngineVGA_reset),
    .io_spriteXPosition_0(graphicEngineVGA_io_spriteXPosition_0),
    .io_spriteXPosition_1(graphicEngineVGA_io_spriteXPosition_1),
    .io_spriteXPosition_2(graphicEngineVGA_io_spriteXPosition_2),
    .io_spriteXPosition_3(graphicEngineVGA_io_spriteXPosition_3),
    .io_spriteXPosition_4(graphicEngineVGA_io_spriteXPosition_4),
    .io_spriteXPosition_5(graphicEngineVGA_io_spriteXPosition_5),
    .io_spriteXPosition_6(graphicEngineVGA_io_spriteXPosition_6),
    .io_spriteXPosition_7(graphicEngineVGA_io_spriteXPosition_7),
    .io_spriteXPosition_8(graphicEngineVGA_io_spriteXPosition_8),
    .io_spriteXPosition_9(graphicEngineVGA_io_spriteXPosition_9),
    .io_spriteXPosition_10(graphicEngineVGA_io_spriteXPosition_10),
    .io_spriteXPosition_11(graphicEngineVGA_io_spriteXPosition_11),
    .io_spriteXPosition_12(graphicEngineVGA_io_spriteXPosition_12),
    .io_spriteXPosition_13(graphicEngineVGA_io_spriteXPosition_13),
    .io_spriteXPosition_14(graphicEngineVGA_io_spriteXPosition_14),
    .io_spriteXPosition_15(graphicEngineVGA_io_spriteXPosition_15),
    .io_spriteXPosition_16(graphicEngineVGA_io_spriteXPosition_16),
    .io_spriteXPosition_17(graphicEngineVGA_io_spriteXPosition_17),
    .io_spriteXPosition_18(graphicEngineVGA_io_spriteXPosition_18),
    .io_spriteXPosition_19(graphicEngineVGA_io_spriteXPosition_19),
    .io_spriteXPosition_20(graphicEngineVGA_io_spriteXPosition_20),
    .io_spriteXPosition_21(graphicEngineVGA_io_spriteXPosition_21),
    .io_spriteXPosition_22(graphicEngineVGA_io_spriteXPosition_22),
    .io_spriteXPosition_23(graphicEngineVGA_io_spriteXPosition_23),
    .io_spriteXPosition_24(graphicEngineVGA_io_spriteXPosition_24),
    .io_spriteXPosition_25(graphicEngineVGA_io_spriteXPosition_25),
    .io_spriteXPosition_26(graphicEngineVGA_io_spriteXPosition_26),
    .io_spriteXPosition_27(graphicEngineVGA_io_spriteXPosition_27),
    .io_spriteYPosition_0(graphicEngineVGA_io_spriteYPosition_0),
    .io_spriteYPosition_1(graphicEngineVGA_io_spriteYPosition_1),
    .io_spriteYPosition_2(graphicEngineVGA_io_spriteYPosition_2),
    .io_spriteYPosition_3(graphicEngineVGA_io_spriteYPosition_3),
    .io_spriteYPosition_4(graphicEngineVGA_io_spriteYPosition_4),
    .io_spriteYPosition_5(graphicEngineVGA_io_spriteYPosition_5),
    .io_spriteYPosition_6(graphicEngineVGA_io_spriteYPosition_6),
    .io_spriteYPosition_7(graphicEngineVGA_io_spriteYPosition_7),
    .io_spriteYPosition_8(graphicEngineVGA_io_spriteYPosition_8),
    .io_spriteYPosition_9(graphicEngineVGA_io_spriteYPosition_9),
    .io_spriteYPosition_10(graphicEngineVGA_io_spriteYPosition_10),
    .io_spriteYPosition_11(graphicEngineVGA_io_spriteYPosition_11),
    .io_spriteYPosition_12(graphicEngineVGA_io_spriteYPosition_12),
    .io_spriteYPosition_13(graphicEngineVGA_io_spriteYPosition_13),
    .io_spriteYPosition_14(graphicEngineVGA_io_spriteYPosition_14),
    .io_spriteYPosition_15(graphicEngineVGA_io_spriteYPosition_15),
    .io_spriteYPosition_16(graphicEngineVGA_io_spriteYPosition_16),
    .io_spriteYPosition_17(graphicEngineVGA_io_spriteYPosition_17),
    .io_spriteYPosition_18(graphicEngineVGA_io_spriteYPosition_18),
    .io_spriteYPosition_19(graphicEngineVGA_io_spriteYPosition_19),
    .io_spriteYPosition_20(graphicEngineVGA_io_spriteYPosition_20),
    .io_spriteYPosition_21(graphicEngineVGA_io_spriteYPosition_21),
    .io_spriteYPosition_22(graphicEngineVGA_io_spriteYPosition_22),
    .io_spriteYPosition_23(graphicEngineVGA_io_spriteYPosition_23),
    .io_spriteYPosition_24(graphicEngineVGA_io_spriteYPosition_24),
    .io_spriteYPosition_25(graphicEngineVGA_io_spriteYPosition_25),
    .io_spriteYPosition_26(graphicEngineVGA_io_spriteYPosition_26),
    .io_spriteYPosition_27(graphicEngineVGA_io_spriteYPosition_27),
    .io_spriteVisible_0(graphicEngineVGA_io_spriteVisible_0),
    .io_spriteVisible_1(graphicEngineVGA_io_spriteVisible_1),
    .io_spriteVisible_2(graphicEngineVGA_io_spriteVisible_2),
    .io_spriteVisible_3(graphicEngineVGA_io_spriteVisible_3),
    .io_spriteVisible_4(graphicEngineVGA_io_spriteVisible_4),
    .io_spriteVisible_5(graphicEngineVGA_io_spriteVisible_5),
    .io_spriteVisible_6(graphicEngineVGA_io_spriteVisible_6),
    .io_spriteVisible_7(graphicEngineVGA_io_spriteVisible_7),
    .io_spriteVisible_8(graphicEngineVGA_io_spriteVisible_8),
    .io_spriteVisible_9(graphicEngineVGA_io_spriteVisible_9),
    .io_spriteVisible_10(graphicEngineVGA_io_spriteVisible_10),
    .io_spriteVisible_11(graphicEngineVGA_io_spriteVisible_11),
    .io_spriteVisible_12(graphicEngineVGA_io_spriteVisible_12),
    .io_spriteVisible_13(graphicEngineVGA_io_spriteVisible_13),
    .io_spriteVisible_14(graphicEngineVGA_io_spriteVisible_14),
    .io_spriteVisible_15(graphicEngineVGA_io_spriteVisible_15),
    .io_spriteVisible_16(graphicEngineVGA_io_spriteVisible_16),
    .io_spriteVisible_17(graphicEngineVGA_io_spriteVisible_17),
    .io_spriteVisible_18(graphicEngineVGA_io_spriteVisible_18),
    .io_spriteVisible_19(graphicEngineVGA_io_spriteVisible_19),
    .io_spriteVisible_20(graphicEngineVGA_io_spriteVisible_20),
    .io_spriteVisible_21(graphicEngineVGA_io_spriteVisible_21),
    .io_spriteVisible_22(graphicEngineVGA_io_spriteVisible_22),
    .io_spriteVisible_23(graphicEngineVGA_io_spriteVisible_23),
    .io_spriteVisible_24(graphicEngineVGA_io_spriteVisible_24),
    .io_spriteVisible_25(graphicEngineVGA_io_spriteVisible_25),
    .io_spriteVisible_26(graphicEngineVGA_io_spriteVisible_26),
    .io_spriteVisible_27(graphicEngineVGA_io_spriteVisible_27),
    .io_viewBoxX(graphicEngineVGA_io_viewBoxX),
    .io_viewBoxY(graphicEngineVGA_io_viewBoxY),
    .io_backBufferWriteData(graphicEngineVGA_io_backBufferWriteData),
    .io_backBufferWriteAddress(graphicEngineVGA_io_backBufferWriteAddress),
    .io_backBufferWriteEnable(graphicEngineVGA_io_backBufferWriteEnable),
    .io_newFrame(graphicEngineVGA_io_newFrame),
    .io_frameUpdateDone(graphicEngineVGA_io_frameUpdateDone),
    .io_missingFrameError(graphicEngineVGA_io_missingFrameError),
    .io_backBufferWriteError(graphicEngineVGA_io_backBufferWriteError),
    .io_viewBoxOutOfRangeError(graphicEngineVGA_io_viewBoxOutOfRangeError),
    .io_vgaRed(graphicEngineVGA_io_vgaRed),
    .io_vgaBlue(graphicEngineVGA_io_vgaBlue),
    .io_vgaGreen(graphicEngineVGA_io_vgaGreen),
    .io_Hsync(graphicEngineVGA_io_Hsync),
    .io_Vsync(graphicEngineVGA_io_Vsync)
  );
  SoundEngine soundEngine ( // @[\\src\\main\\scala\\GameTop.scala 49:27]
    .clock(soundEngine_clock),
    .reset(soundEngine_reset),
    .io_soundOut(soundEngine_io_soundOut),
    .io_startTune_0(soundEngine_io_startTune_0)
  );
  GameLogic gameLogic ( // @[\\src\\main\\scala\\GameTop.scala 53:25]
    .clock(gameLogic_clock),
    .reset(gameLogic_reset),
    .io_btnU(gameLogic_io_btnU),
    .io_btnL(gameLogic_io_btnL),
    .io_btnR(gameLogic_io_btnR),
    .io_btnD(gameLogic_io_btnD),
    .io_sw_7(gameLogic_io_sw_7),
    .io_led_0(gameLogic_io_led_0),
    .io_led_1(gameLogic_io_led_1),
    .io_led_2(gameLogic_io_led_2),
    .io_led_3(gameLogic_io_led_3),
    .io_spriteXPosition_0(gameLogic_io_spriteXPosition_0),
    .io_spriteXPosition_1(gameLogic_io_spriteXPosition_1),
    .io_spriteXPosition_2(gameLogic_io_spriteXPosition_2),
    .io_spriteXPosition_3(gameLogic_io_spriteXPosition_3),
    .io_spriteXPosition_4(gameLogic_io_spriteXPosition_4),
    .io_spriteXPosition_5(gameLogic_io_spriteXPosition_5),
    .io_spriteXPosition_6(gameLogic_io_spriteXPosition_6),
    .io_spriteXPosition_7(gameLogic_io_spriteXPosition_7),
    .io_spriteXPosition_8(gameLogic_io_spriteXPosition_8),
    .io_spriteXPosition_9(gameLogic_io_spriteXPosition_9),
    .io_spriteXPosition_10(gameLogic_io_spriteXPosition_10),
    .io_spriteXPosition_11(gameLogic_io_spriteXPosition_11),
    .io_spriteXPosition_12(gameLogic_io_spriteXPosition_12),
    .io_spriteXPosition_13(gameLogic_io_spriteXPosition_13),
    .io_spriteXPosition_14(gameLogic_io_spriteXPosition_14),
    .io_spriteXPosition_15(gameLogic_io_spriteXPosition_15),
    .io_spriteXPosition_16(gameLogic_io_spriteXPosition_16),
    .io_spriteXPosition_17(gameLogic_io_spriteXPosition_17),
    .io_spriteXPosition_18(gameLogic_io_spriteXPosition_18),
    .io_spriteXPosition_19(gameLogic_io_spriteXPosition_19),
    .io_spriteXPosition_20(gameLogic_io_spriteXPosition_20),
    .io_spriteXPosition_21(gameLogic_io_spriteXPosition_21),
    .io_spriteXPosition_22(gameLogic_io_spriteXPosition_22),
    .io_spriteXPosition_23(gameLogic_io_spriteXPosition_23),
    .io_spriteXPosition_24(gameLogic_io_spriteXPosition_24),
    .io_spriteXPosition_25(gameLogic_io_spriteXPosition_25),
    .io_spriteXPosition_26(gameLogic_io_spriteXPosition_26),
    .io_spriteXPosition_27(gameLogic_io_spriteXPosition_27),
    .io_spriteYPosition_0(gameLogic_io_spriteYPosition_0),
    .io_spriteYPosition_1(gameLogic_io_spriteYPosition_1),
    .io_spriteYPosition_2(gameLogic_io_spriteYPosition_2),
    .io_spriteYPosition_3(gameLogic_io_spriteYPosition_3),
    .io_spriteYPosition_4(gameLogic_io_spriteYPosition_4),
    .io_spriteYPosition_5(gameLogic_io_spriteYPosition_5),
    .io_spriteYPosition_6(gameLogic_io_spriteYPosition_6),
    .io_spriteYPosition_7(gameLogic_io_spriteYPosition_7),
    .io_spriteYPosition_8(gameLogic_io_spriteYPosition_8),
    .io_spriteYPosition_9(gameLogic_io_spriteYPosition_9),
    .io_spriteYPosition_10(gameLogic_io_spriteYPosition_10),
    .io_spriteYPosition_11(gameLogic_io_spriteYPosition_11),
    .io_spriteYPosition_12(gameLogic_io_spriteYPosition_12),
    .io_spriteYPosition_13(gameLogic_io_spriteYPosition_13),
    .io_spriteYPosition_14(gameLogic_io_spriteYPosition_14),
    .io_spriteYPosition_15(gameLogic_io_spriteYPosition_15),
    .io_spriteYPosition_16(gameLogic_io_spriteYPosition_16),
    .io_spriteYPosition_17(gameLogic_io_spriteYPosition_17),
    .io_spriteYPosition_18(gameLogic_io_spriteYPosition_18),
    .io_spriteYPosition_19(gameLogic_io_spriteYPosition_19),
    .io_spriteYPosition_20(gameLogic_io_spriteYPosition_20),
    .io_spriteYPosition_21(gameLogic_io_spriteYPosition_21),
    .io_spriteYPosition_22(gameLogic_io_spriteYPosition_22),
    .io_spriteYPosition_23(gameLogic_io_spriteYPosition_23),
    .io_spriteYPosition_24(gameLogic_io_spriteYPosition_24),
    .io_spriteYPosition_25(gameLogic_io_spriteYPosition_25),
    .io_spriteYPosition_26(gameLogic_io_spriteYPosition_26),
    .io_spriteYPosition_27(gameLogic_io_spriteYPosition_27),
    .io_spriteVisible_0(gameLogic_io_spriteVisible_0),
    .io_spriteVisible_1(gameLogic_io_spriteVisible_1),
    .io_spriteVisible_2(gameLogic_io_spriteVisible_2),
    .io_spriteVisible_3(gameLogic_io_spriteVisible_3),
    .io_spriteVisible_4(gameLogic_io_spriteVisible_4),
    .io_spriteVisible_5(gameLogic_io_spriteVisible_5),
    .io_spriteVisible_6(gameLogic_io_spriteVisible_6),
    .io_spriteVisible_7(gameLogic_io_spriteVisible_7),
    .io_spriteVisible_8(gameLogic_io_spriteVisible_8),
    .io_spriteVisible_9(gameLogic_io_spriteVisible_9),
    .io_spriteVisible_10(gameLogic_io_spriteVisible_10),
    .io_spriteVisible_11(gameLogic_io_spriteVisible_11),
    .io_spriteVisible_12(gameLogic_io_spriteVisible_12),
    .io_spriteVisible_13(gameLogic_io_spriteVisible_13),
    .io_spriteVisible_14(gameLogic_io_spriteVisible_14),
    .io_spriteVisible_15(gameLogic_io_spriteVisible_15),
    .io_spriteVisible_16(gameLogic_io_spriteVisible_16),
    .io_spriteVisible_17(gameLogic_io_spriteVisible_17),
    .io_spriteVisible_18(gameLogic_io_spriteVisible_18),
    .io_spriteVisible_19(gameLogic_io_spriteVisible_19),
    .io_spriteVisible_20(gameLogic_io_spriteVisible_20),
    .io_spriteVisible_21(gameLogic_io_spriteVisible_21),
    .io_spriteVisible_22(gameLogic_io_spriteVisible_22),
    .io_spriteVisible_23(gameLogic_io_spriteVisible_23),
    .io_spriteVisible_24(gameLogic_io_spriteVisible_24),
    .io_spriteVisible_25(gameLogic_io_spriteVisible_25),
    .io_spriteVisible_26(gameLogic_io_spriteVisible_26),
    .io_spriteVisible_27(gameLogic_io_spriteVisible_27),
    .io_viewBoxX(gameLogic_io_viewBoxX),
    .io_viewBoxY(gameLogic_io_viewBoxY),
    .io_backBufferWriteData(gameLogic_io_backBufferWriteData),
    .io_backBufferWriteAddress(gameLogic_io_backBufferWriteAddress),
    .io_backBufferWriteEnable(gameLogic_io_backBufferWriteEnable),
    .io_newFrame(gameLogic_io_newFrame),
    .io_frameUpdateDone(gameLogic_io_frameUpdateDone),
    .io_startTune_0(gameLogic_io_startTune_0)
  );
  assign io_vgaRed = graphicEngineVGA_io_vgaRed; // @[\\src\\main\\scala\\GameTop.scala 96:13]
  assign io_vgaBlue = graphicEngineVGA_io_vgaBlue; // @[\\src\\main\\scala\\GameTop.scala 98:14]
  assign io_vgaGreen = graphicEngineVGA_io_vgaGreen; // @[\\src\\main\\scala\\GameTop.scala 97:15]
  assign io_Hsync = graphicEngineVGA_io_Hsync; // @[\\src\\main\\scala\\GameTop.scala 99:12]
  assign io_Vsync = graphicEngineVGA_io_Vsync; // @[\\src\\main\\scala\\GameTop.scala 100:12]
  assign io_led_0 = gameLogic_io_led_0; // @[\\src\\main\\scala\\GameTop.scala 108:10]
  assign io_led_1 = gameLogic_io_led_1; // @[\\src\\main\\scala\\GameTop.scala 108:10]
  assign io_led_2 = gameLogic_io_led_2; // @[\\src\\main\\scala\\GameTop.scala 108:10]
  assign io_led_3 = gameLogic_io_led_3; // @[\\src\\main\\scala\\GameTop.scala 108:10]
  assign io_missingFrameError = graphicEngineVGA_io_missingFrameError; // @[\\src\\main\\scala\\GameTop.scala 111:24]
  assign io_backBufferWriteError = graphicEngineVGA_io_backBufferWriteError; // @[\\src\\main\\scala\\GameTop.scala 112:27]
  assign io_viewBoxOutOfRangeError = graphicEngineVGA_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\GameTop.scala 113:29]
  assign io_soundOut = soundEngine_io_soundOut; // @[\\src\\main\\scala\\GameTop.scala 142:15]
  assign graphicEngineVGA_clock = clock;
  assign graphicEngineVGA_reset = resetReleaseCounter == 22'h3d08ff ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameTop.scala 74:67 75:18 77:18]
  assign graphicEngineVGA_io_spriteXPosition_0 = gameLogic_io_spriteXPosition_0; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_1 = gameLogic_io_spriteXPosition_1; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_2 = gameLogic_io_spriteXPosition_2; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_3 = gameLogic_io_spriteXPosition_3; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_4 = gameLogic_io_spriteXPosition_4; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_5 = gameLogic_io_spriteXPosition_5; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_6 = gameLogic_io_spriteXPosition_6; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_7 = gameLogic_io_spriteXPosition_7; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_8 = gameLogic_io_spriteXPosition_8; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_9 = gameLogic_io_spriteXPosition_9; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_10 = gameLogic_io_spriteXPosition_10; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_11 = gameLogic_io_spriteXPosition_11; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_12 = gameLogic_io_spriteXPosition_12; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_13 = gameLogic_io_spriteXPosition_13; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_14 = gameLogic_io_spriteXPosition_14; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_15 = gameLogic_io_spriteXPosition_15; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_16 = gameLogic_io_spriteXPosition_16; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_17 = gameLogic_io_spriteXPosition_17; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_18 = gameLogic_io_spriteXPosition_18; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_19 = gameLogic_io_spriteXPosition_19; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_20 = gameLogic_io_spriteXPosition_20; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_21 = gameLogic_io_spriteXPosition_21; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_22 = gameLogic_io_spriteXPosition_22; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_23 = gameLogic_io_spriteXPosition_23; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_24 = gameLogic_io_spriteXPosition_24; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_25 = gameLogic_io_spriteXPosition_25; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_26 = gameLogic_io_spriteXPosition_26; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteXPosition_27 = gameLogic_io_spriteXPosition_27; // @[\\src\\main\\scala\\GameTop.scala 116:39]
  assign graphicEngineVGA_io_spriteYPosition_0 = gameLogic_io_spriteYPosition_0; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_1 = gameLogic_io_spriteYPosition_1; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_2 = gameLogic_io_spriteYPosition_2; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_3 = gameLogic_io_spriteYPosition_3; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_4 = gameLogic_io_spriteYPosition_4; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_5 = gameLogic_io_spriteYPosition_5; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_6 = gameLogic_io_spriteYPosition_6; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_7 = gameLogic_io_spriteYPosition_7; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_8 = gameLogic_io_spriteYPosition_8; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_9 = gameLogic_io_spriteYPosition_9; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_10 = gameLogic_io_spriteYPosition_10; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_11 = gameLogic_io_spriteYPosition_11; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_12 = gameLogic_io_spriteYPosition_12; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_13 = gameLogic_io_spriteYPosition_13; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_14 = gameLogic_io_spriteYPosition_14; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_15 = gameLogic_io_spriteYPosition_15; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_16 = gameLogic_io_spriteYPosition_16; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_17 = gameLogic_io_spriteYPosition_17; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_18 = gameLogic_io_spriteYPosition_18; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_19 = gameLogic_io_spriteYPosition_19; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_20 = gameLogic_io_spriteYPosition_20; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_21 = gameLogic_io_spriteYPosition_21; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_22 = gameLogic_io_spriteYPosition_22; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_23 = gameLogic_io_spriteYPosition_23; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_24 = gameLogic_io_spriteYPosition_24; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_25 = gameLogic_io_spriteYPosition_25; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_26 = gameLogic_io_spriteYPosition_26; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteYPosition_27 = gameLogic_io_spriteYPosition_27; // @[\\src\\main\\scala\\GameTop.scala 117:39]
  assign graphicEngineVGA_io_spriteVisible_0 = gameLogic_io_spriteVisible_0; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_1 = gameLogic_io_spriteVisible_1; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_2 = gameLogic_io_spriteVisible_2; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_3 = gameLogic_io_spriteVisible_3; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_4 = gameLogic_io_spriteVisible_4; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_5 = gameLogic_io_spriteVisible_5; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_6 = gameLogic_io_spriteVisible_6; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_7 = gameLogic_io_spriteVisible_7; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_8 = gameLogic_io_spriteVisible_8; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_9 = gameLogic_io_spriteVisible_9; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_10 = gameLogic_io_spriteVisible_10; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_11 = gameLogic_io_spriteVisible_11; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_12 = gameLogic_io_spriteVisible_12; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_13 = gameLogic_io_spriteVisible_13; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_14 = gameLogic_io_spriteVisible_14; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_15 = gameLogic_io_spriteVisible_15; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_16 = gameLogic_io_spriteVisible_16; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_17 = gameLogic_io_spriteVisible_17; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_18 = gameLogic_io_spriteVisible_18; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_19 = gameLogic_io_spriteVisible_19; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_20 = gameLogic_io_spriteVisible_20; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_21 = gameLogic_io_spriteVisible_21; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_22 = gameLogic_io_spriteVisible_22; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_23 = gameLogic_io_spriteVisible_23; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_24 = gameLogic_io_spriteVisible_24; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_25 = gameLogic_io_spriteVisible_25; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_26 = gameLogic_io_spriteVisible_26; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_spriteVisible_27 = gameLogic_io_spriteVisible_27; // @[\\src\\main\\scala\\GameTop.scala 118:37]
  assign graphicEngineVGA_io_viewBoxX = gameLogic_io_viewBoxX; // @[\\src\\main\\scala\\GameTop.scala 129:32]
  assign graphicEngineVGA_io_viewBoxY = gameLogic_io_viewBoxY; // @[\\src\\main\\scala\\GameTop.scala 130:32]
  assign graphicEngineVGA_io_backBufferWriteData = gameLogic_io_backBufferWriteData; // @[\\src\\main\\scala\\GameTop.scala 133:43]
  assign graphicEngineVGA_io_backBufferWriteAddress = gameLogic_io_backBufferWriteAddress; // @[\\src\\main\\scala\\GameTop.scala 134:46]
  assign graphicEngineVGA_io_backBufferWriteEnable = gameLogic_io_backBufferWriteEnable; // @[\\src\\main\\scala\\GameTop.scala 135:45]
  assign graphicEngineVGA_io_frameUpdateDone = gameLogic_io_frameUpdateDone; // @[\\src\\main\\scala\\GameTop.scala 139:39]
  assign soundEngine_clock = clock;
  assign soundEngine_reset = reset;
  assign soundEngine_io_startTune_0 = gameLogic_io_startTune_0; // @[\\src\\main\\scala\\GameTop.scala 143:28]
  assign gameLogic_clock = clock;
  assign gameLogic_reset = resetReleaseCounter == 22'h3d08ff ? 1'h0 : 1'h1; // @[\\src\\main\\scala\\GameTop.scala 74:67 75:18 77:18]
  assign gameLogic_io_btnU = btnUState; // @[\\src\\main\\scala\\GameTop.scala 90:21]
  assign gameLogic_io_btnL = btnLState; // @[\\src\\main\\scala\\GameTop.scala 91:21]
  assign gameLogic_io_btnR = btnRState; // @[\\src\\main\\scala\\GameTop.scala 92:21]
  assign gameLogic_io_btnD = btnDState; // @[\\src\\main\\scala\\GameTop.scala 93:21]
  assign gameLogic_io_sw_7 = gameLogic_io_sw_7_r; // @[\\src\\main\\scala\\GameTop.scala 104:24]
  assign gameLogic_io_newFrame = graphicEngineVGA_io_newFrame; // @[\\src\\main\\scala\\GameTop.scala 138:25]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 59:32]
      debounceCounter <= 21'h0; // @[\\src\\main\\scala\\GameTop.scala 59:32]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 61:57]
      debounceCounter <= 21'h0; // @[\\src\\main\\scala\\GameTop.scala 62:21]
    end else begin
      debounceCounter <= _debounceCounter_T_1; // @[\\src\\main\\scala\\GameTop.scala 65:21]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 72:36]
      resetReleaseCounter <= 22'h0; // @[\\src\\main\\scala\\GameTop.scala 72:36]
    end else if (!(resetReleaseCounter == 22'h3d08ff)) begin // @[\\src\\main\\scala\\GameTop.scala 74:67]
      resetReleaseCounter <= _resetReleaseCounter_T_1; // @[\\src\\main\\scala\\GameTop.scala 78:25]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_0 <= btnUState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_1 <= btnUState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnUState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnUState_pipeReg_2 <= io_btnU; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 85:28]
      btnUState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 85:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 85:28]
      btnUState <= btnUState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 85:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_0 <= btnLState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_1 <= btnLState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnLState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnLState_pipeReg_2 <= io_btnL; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 86:28]
      btnLState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 86:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 86:28]
      btnLState <= btnLState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 86:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_0 <= btnRState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_1 <= btnRState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnRState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnRState_pipeReg_2 <= io_btnR; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 87:28]
      btnRState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 87:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 87:28]
      btnRState <= btnRState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 87:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_0 <= btnDState_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_1 <= btnDState_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      btnDState_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      btnDState_pipeReg_2 <= io_btnD; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 88:28]
      btnDState <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 88:28]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 88:28]
      btnDState <= btnDState_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 88:28]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      gameLogic_io_sw_7_pipeReg_0 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      gameLogic_io_sw_7_pipeReg_0 <= gameLogic_io_sw_7_pipeReg_1; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      gameLogic_io_sw_7_pipeReg_1 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      gameLogic_io_sw_7_pipeReg_1 <= gameLogic_io_sw_7_pipeReg_2; // @[\\src\\main\\scala\\GameUtilities.scala 43:20]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
      gameLogic_io_sw_7_pipeReg_2 <= 1'h0; // @[\\src\\main\\scala\\GameUtilities.scala 39:28]
    end else begin
      gameLogic_io_sw_7_pipeReg_2 <= io_sw_7; // @[\\src\\main\\scala\\GameUtilities.scala 41:30]
    end
    if (reset) begin // @[\\src\\main\\scala\\GameTop.scala 104:36]
      gameLogic_io_sw_7_r <= 1'h0; // @[\\src\\main\\scala\\GameTop.scala 104:36]
    end else if (debounceSampleEn) begin // @[\\src\\main\\scala\\GameTop.scala 104:36]
      gameLogic_io_sw_7_r <= gameLogic_io_sw_7_pipeReg_0; // @[\\src\\main\\scala\\GameTop.scala 104:36]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounceCounter = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  resetReleaseCounter = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btnUState_pipeReg_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  btnUState_pipeReg_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  btnUState_pipeReg_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  btnUState = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  btnLState_pipeReg_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  btnLState_pipeReg_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  btnLState_pipeReg_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btnLState = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  btnRState_pipeReg_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  btnRState_pipeReg_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  btnRState_pipeReg_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btnRState = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  btnDState_pipeReg_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  btnDState_pipeReg_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  btnDState_pipeReg_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  btnDState = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  gameLogic_io_sw_7_pipeReg_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  gameLogic_io_sw_7_pipeReg_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  gameLogic_io_sw_7_pipeReg_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  gameLogic_io_sw_7_r = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input        clock,
  input        reset,
  input        io_btnC, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnU, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnL, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnR, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_btnD, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaRed, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaGreen, // @[\\src\\main\\scala\\Top.scala 14:14]
  output [3:0] io_vgaBlue, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_Hsync, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_Vsync, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_0, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_1, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_2, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_3, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_4, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_5, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_6, // @[\\src\\main\\scala\\Top.scala 14:14]
  input        io_sw_7, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_0, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_1, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_2, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_3, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_4, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_5, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_6, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_led_7, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_missingFrameError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_backBufferWriteError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_viewBoxOutOfRangeError, // @[\\src\\main\\scala\\Top.scala 14:14]
  output       io_soundOut // @[\\src\\main\\scala\\Top.scala 14:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  gameTop_clock; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_reset; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnU; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnL; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnR; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_btnD; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaRed; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaBlue; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire [3:0] gameTop_io_vgaGreen; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_Hsync; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_Vsync; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_sw_7; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_led_0; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_led_1; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_led_2; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_led_3; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_missingFrameError; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_backBufferWriteError; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\Top.scala 44:23]
  wire  gameTop_io_soundOut; // @[\\src\\main\\scala\\Top.scala 44:23]
  reg  syncResetInput_REG; // @[\\src\\main\\scala\\Top.scala 49:48]
  reg  syncResetInput_REG_1; // @[\\src\\main\\scala\\Top.scala 49:40]
  reg  syncResetInput_REG_2; // @[\\src\\main\\scala\\Top.scala 49:32]
  reg  pipeResetReg_0; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_1; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_2; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_3; // @[\\src\\main\\scala\\Top.scala 54:25]
  reg  pipeResetReg_4; // @[\\src\\main\\scala\\Top.scala 54:25]
  wire [4:0] _gameTop_reset_T = {pipeResetReg_4,pipeResetReg_3,pipeResetReg_2,pipeResetReg_1,pipeResetReg_0}; // @[\\src\\main\\scala\\Top.scala 59:33]
  GameTop gameTop ( // @[\\src\\main\\scala\\Top.scala 44:23]
    .clock(gameTop_clock),
    .reset(gameTop_reset),
    .io_btnU(gameTop_io_btnU),
    .io_btnL(gameTop_io_btnL),
    .io_btnR(gameTop_io_btnR),
    .io_btnD(gameTop_io_btnD),
    .io_vgaRed(gameTop_io_vgaRed),
    .io_vgaBlue(gameTop_io_vgaBlue),
    .io_vgaGreen(gameTop_io_vgaGreen),
    .io_Hsync(gameTop_io_Hsync),
    .io_Vsync(gameTop_io_Vsync),
    .io_sw_7(gameTop_io_sw_7),
    .io_led_0(gameTop_io_led_0),
    .io_led_1(gameTop_io_led_1),
    .io_led_2(gameTop_io_led_2),
    .io_led_3(gameTop_io_led_3),
    .io_missingFrameError(gameTop_io_missingFrameError),
    .io_backBufferWriteError(gameTop_io_backBufferWriteError),
    .io_viewBoxOutOfRangeError(gameTop_io_viewBoxOutOfRangeError),
    .io_soundOut(gameTop_io_soundOut)
  );
  assign io_vgaRed = gameTop_io_vgaRed; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_vgaGreen = gameTop_io_vgaGreen; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_vgaBlue = gameTop_io_vgaBlue; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_Hsync = gameTop_io_Hsync; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_Vsync = gameTop_io_Vsync; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_0 = gameTop_io_led_0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_1 = gameTop_io_led_1; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_2 = gameTop_io_led_2; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_3 = gameTop_io_led_3; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_4 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_5 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_6 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_led_7 = 1'h0; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_missingFrameError = gameTop_io_missingFrameError; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_backBufferWriteError = gameTop_io_backBufferWriteError; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_viewBoxOutOfRangeError = gameTop_io_viewBoxOutOfRangeError; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign io_soundOut = gameTop_io_soundOut; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_clock = clock;
  assign gameTop_reset = |_gameTop_reset_T; // @[\\src\\main\\scala\\Top.scala 59:40]
  assign gameTop_io_btnU = io_btnU; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnL = io_btnL; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnR = io_btnR; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_btnD = io_btnD; // @[\\src\\main\\scala\\Top.scala 62:14]
  assign gameTop_io_sw_7 = io_sw_7; // @[\\src\\main\\scala\\Top.scala 62:14]
  always @(posedge clock) begin
    syncResetInput_REG <= reset; // @[\\src\\main\\scala\\Top.scala 49:48]
    syncResetInput_REG_1 <= syncResetInput_REG; // @[\\src\\main\\scala\\Top.scala 49:40]
    syncResetInput_REG_2 <= syncResetInput_REG_1; // @[\\src\\main\\scala\\Top.scala 49:32]
    pipeResetReg_0 <= pipeResetReg_1; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_1 <= pipeResetReg_2; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_2 <= pipeResetReg_3; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_3 <= pipeResetReg_4; // @[\\src\\main\\scala\\Top.scala 57:21]
    pipeResetReg_4 <= ~syncResetInput_REG_2; // @[\\src\\main\\scala\\Top.scala 49:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  syncResetInput_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  syncResetInput_REG_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  syncResetInput_REG_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pipeResetReg_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pipeResetReg_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pipeResetReg_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pipeResetReg_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pipeResetReg_4 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
